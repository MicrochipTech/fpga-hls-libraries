--=================================================================================================
-- File Name                           : VGA_Controller_SHLS.vhd
-- Description                         : Supporting both Native mode and AXI4 Stream mode
-- Targeted device                     : Microsemi-SoC
-- Author                              : India Solutions Team
--
-- COPYRIGHT 2021 BY MICROSEMI
-- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS FROM MICROSEMI
-- CORP. IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM MICROSEMI FOR USE OF THIS
-- FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND NO BACK-UP OF THE FILE SHOULD BE MADE.
--
--=================================================================================================
--=================================================================================================
-- Libraries
--=================================================================================================
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
--=================================================================================================
-- VGA_Controller_SHLS entity declaration
--=================================================================================================                                                                                                                          
entity VGA_Controller_SHLS is
  generic(
-- Generic List
    -- Video format selection
    g_VIDEO_FORMAT : integer := 1;  -- 0 -> 1280x720 1 -> 1920x1080 2-> 3840x2160 3-> 640x360

    g_PIXELS_PER_CLK : integer := 1;

    G_FORMAT : integer := 0;  --  0= VGA_Controller_SHLS and 1= VGA_Controller_SHLS with AXI       

    --Added for AXIS_Video
    g_FIFO_WIDTHAD :integer := 3 -- FIFO address width
    );
  port (
-- Port List
    -------------------------------------------------------------------------------------------------------------------------------
    --Added for AXIS_Video
    --begin
    --start of frame
    SOF : in std_logic;

    --End of line
    EOL : in std_logic;

    --Pop FIFO (used to pop FIFO during the alignment phase)
    POP_FIFO : out std_logic;

    --number of words in FIFO
    FIFO_FILL_LVL : in std_logic_vector(g_FIFO_WIDTHAD downto 0);

    --FIFO almost empty
    FIFO_AE : in std_logic;

    --AXI Tvalid
    AXI_VALID : in std_logic;

   
    --end
    ------------------------------------------------------------------------------------------------------------------------------
    
    -- System reset
    RESETN_I : in std_logic;

    -- System clock
    SYS_CLK_I : in std_logic;

    -- Specifies enable
    ENABLE_I : in std_logic;

    -- enable external syncing
    ENABLE_EXT_SYNC_I : in std_logic;

    -- external sync reference signal
    -- EXT_SYNC_SIGNAL_I : in std_logic;

    -- Specifies the valid control signal
    TVALID_I : in std_logic;

    TREADY_O : out std_logic;
    -- Active horizontal sync pulse
    H_SYNC_O : out std_logic;

    -- Active vertical sync pulse
    V_SYNC_O : out std_logic;

    -- Data trigger
    DATA_TRIGGER_O : out std_logic;

    -- Frame end
    FRAME_END_O : out std_logic;

    -- Data Enable
    DATA_ENABLE_O : out std_logic;

    -- Display data (used to indicate video data is stable so incoming data will be displayed instead of yellow screen)
    DISPLAY_DATA_O : out std_logic;


    V_ACTIVE_O : out std_logic;

    --Horizontal Resolution
    H_RES_O : out std_logic_vector(15 downto 0);

    TDATA_O : out std_logic_vector(7 downto 0);

    TSTRB_O : out std_logic_vector(2 downto 0);

    TKEEP_O : out std_logic_vector(2 downto 0);
    TUSER_O : out std_logic_vector(3 downto 0);

    TLAST_O : out std_logic;

    -- Specifies the valid control signal
    TVALID_O : out std_logic

    );
end VGA_Controller_SHLS;

`protect begin_protected
`protect version=1
`protect author="Alireza Mellat", author_info="Software Engineer - Microchip"
`protect encrypt_agent="encryptP1735.pl", encrypt_agent_info="Synplify encryption scripts"

`protect key_keyowner="Synplicity", key_keyname="SYNP05_001", key_method="rsa"
`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_block
lUI5HtleSvkhs5KELgAkYm3EVy+WVSf9nTAok+qPfZxTUrx4L8WWwHDyJj6rYyInR93txadK4XRy
/Ia08X+YO318Z5lQtcpqRwLSbghn0IhP9IfiT5Q+qVZVUpt8E/X5XZDBsKE0L0zID1NxCNMWLJD/
6VpKIWKLVo8oObY2kjKXlb88y3HAxEiiWC1g3tX3GWKPlh9pm7c3D7a8n9x14o9fMTb5mzTr5mNy
DSBTOV6lJzjE8L+x07MEkUdCezeoTkDvU46q8e8FFUsO0loKPIanjN/z8OUwhnUJUoTVvFcTgqXJ
/5WxhoqtwlOnchDkTPgF0tlsGMXdCaYyyNW4hw==

`protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`protect encoding=(enctype="base64", line_length=76, bytes=128)
`protect key_block
ohZfM36VBAdtp2LteEplqiP0+KOah0NTOf2bEmoSEJv+uy2AQKTWAoIfnP2AFTQz2SOcmHbnHPRN
2XZkNZDx7m/kiMfpJMVr/lAuBSm8xmG4SRuq0yQ14ej1dbhA+8CijMBZ/mFIYMslSMx+14dAzKNv
vvCebdRn7xd4FAUoiIs=

`protect key_keyowner="Microsemi Corporation", key_keyname="MSC-IP-KEY-RSA", key_method="rsa"
`protect encoding=(enctype="base64", line_length=76, bytes=960)
`protect key_block
dP+G7kfagJYQsGMrBG5jbDtMf5PKu9UZwThA2GFiZc4kdQIof4kZMSsItHLhzT7Q9LsIi1VRwo2g
9puiODr1EQ/10aPdSbcsvH75KsWXwP/Nk01QKXSXQjEmbuFMq1rXvfup7C4DkKnzpq5Qnm3wHAoi
cHS43VUVsjrjt4U8a6Bi8nxXJvuAxM14lLL92RiO9t4bBXTvitXoq2DrppsMU+q/X0JV71esxlUJ
Zy86U0hVb88v3KN5FoGtcOYRaGGKXLV6a+wwAWoHznJF+9D9sGGfZCnao7yuJBZxQStQ5TqxiNaR
tFbk2lppj3XzpdSZI/+/XViDL/gssISfzZAmdDOiczytePNttyNFCCxS8vGj1cd8/hI9jGxX3v1D
9x40oo4R2p6vxxSUOP5hb0Wcu4rdABvM2hO2K4wGy2VzI7inh2+n9jYc+QbQP7K1EN7L+TJ2UHuI
wzlrBAJKKTR91ZkGjhBj0RovkNDVrO901FzPTDKPLfi0gt44QtFkKmzjJxayKNHAUm1wphzTuX/I
aGAbAXyH3QtqvL7HucblkkzDRg0+8VH4c4nyeRadzx3XJPPoQJb4A7eapjTBGjUFhCAvq5P/F1UB
tCoOFTZ7cK02jPblZ9IOG5QEZ06urrtd5tzO7uqQdMYH6vQxe17HsjScLH5Ru59IHBPCBgu2gL0v
UE+5Y+4OUzs2fqfTog4qPmdfz+K+XIdFoa3TdEcic6Jg7w+OLFuMWTV01cTn6j86bGXgiBr0hHXD
rGLv3DS21dY4oJIkGvpTsZYh8D3ZhmTR7acyM0lDHJl9dBtTWlQOEof37ipsI1/W1ky0Ep7nqGvA
QEQN3ZXFr0OefmIdb0n/N3KvZ55dUS1ZJBkW/soT073VW83wV+R47GmvM1mKLDG5tGP7IcaHfxQ0
m0QefnyKPzWEQbI4PTnkCghBGLjSoN65vwVQVRZyn38jY69VxDADdB/48EGJj6/kZt+rhFcl1Lq1
YavSg+r/PCsdJDy0K7aHFxVqUnie4ER3wVk/990X7GltnBxjogZtwX1Ep+cgLIGIwSWWbAJlb5nd
OvM1BZnADU9CbuxS2mv8JMwGXBkFumrqrieLZ3yKyNQo2dt7GFV8reAThglwj9JV/FDu7DGm3ttt
4X1kfp2derW/9r1KjZcPMzDTh3jiWozcLnGhDgqWEtPn1CdZa4IOQSTW6yzMp+o8mKff8sHwRXtA
i+FHp+AHYv74YF0DeV5P1vabZtzrTbD1x4Xpp+m1z8QERZC6zTe7TU23vWandT4m

`protect data_keyowner="ip-vendor-a", data_keyname="fpga-ip", data_method="aes128-cbc"
`protect encoding=(enctype="base64", line_length=76, bytes=39168)
`protect data_block
3ilqlGBvNq18mef/zNXgKlK9liUQELfekR6j59np+Dh1fN0RhIN0ZNj/2iJFusUeMJnESHHw8aKW
DQo5ruPvdZSPptmaUOhJ5WpA0joHYIDIgoXlPYD7Aqo5FWkAIhfjlY9oak8dlgNBBBGFf6+cgEws
o0oAh3mz0oBf3upV6Ff1NrCOcRv3mRkIJzpp1J9E6iA8cv/DrZKyHCgstcbNWstuwVD53SPUkGQg
148mwtI+ZF0WqI5IyZjF+JgbyPX2Pj6llmkaq+oCd/r9YDdAWgvIK+6fP5cJtt7rZgSJp65IoVlk
KvGNXBZg1UH/Ko5t2DCB8tt5G5F6IEctaZz3RHkAq5ojOvKR8S00ktxvdgBS5/xThNgUKUi1UiNE
nQxbwu6fon2Mu8/rYA6pzW4KZGovxm0OQX/iajR8mXFcrvosQBUOAdg2g72gerQwouzJbWV0jh8s
dLcPoUk/Uu6xX85fymc408ma/3/WC7ZryWu8EmkMcfhukzJ8u8reTlv9Md5dD4ER/HjCmcj1EpI6
Y7y/USB+S4opkKTW8O+1VKraWZl4+9jMCW8l/TUeuZz0QA5bU54zGX46Xn8ZwvSskeayE1cgkKGt
c9pmzib6C5WSOyiOtVEvSEhiqC8s6g5nLJqT7soQMHDoBsN0Coek4HcQQ3UmD2a8LPRV3R7kWCEn
gyOe3F4dty6EBQ22bmrNqqhfKJzSYD2a65V7AxobBMxRX8d4be14lW2kcDYB2lv55TGlS1yCy8eP
kRM8LzcoFgj4iz4lF0OQLNl+W8VS9fQuqB05WG5C0bWqxxOHY171ppdwviHLI8C6YmWkSyrwnC1l
KYJqqTWx+CoZsjcj7TcGjJFTj5OPLFAK32Rkb6+p9jNYfbrkQ8JHLdh41sXwIgbZzEAz8TEppXKv
0PLBNExK5nAyRWuWOaxuWt9EQeXsDa7+zBBmE1qbww2+TYtFYiI7cM/5Mq/zva5tRv+sAERT6AcY
7pbgvnI6xlMA97i0yPum3TG66BgbXUC2EDZbHeg1U6mot7eBK4gqQpiJ4WemlvWG52+o0HNOR8Jf
maxIbwPosuJpwL0bkLhlZejOB0+1lg7NXwOPRLp/SHapICbx61EtoZkSXoHUXCkJ9/eSo7E6+QK9
D/4uzEMz7av8W9slaqNlPqzQOAa5FYMbSqYo/buuiQyl0Il2XoHeEjz3uNrt1S8RP30zkULug1G+
Hyxfc45Oc5VPSS2ueftx37QznanxY7iP0kxSUS2qDsEY2oiO5EqprxubW2wA4wR/R62fSQzIlPda
GdLeJRZBcJ/r5oBYYFiPSCKFIqARgQmfTnPftV4oxcO7Ygolf40vWJqCmD3lma7smJEDFOmw+DBC
9+6yeaM9tRAJ77hRnnpIEUcxCit5xt3l691WvOROkI8sXUmOVZQiwAHaohFsexThnbT2+fQ62Lda
dvxnf6ODxLuWO+acJ4tnHs4z/j/jhEPRBVzbzCgOM/ztErzdIwifHO/clH2reAM8451/4voXPubi
2G4VWeFCmKzqhxVgd4rrolFTS5PwdKNory54ZQYa6uzQSnmeoea/ovL/HHgmEDKhbWVD0T96OqfV
YB4jm088MlgtjIp+E2IUVgFInnNgn+tklCoR9jgHMcTtDdLfdHQLmB2LhFU1A7cVeIZLYv31UvvK
WDz+xggf62TbGwWp0dJio5v6MpRsgsNyQpbwzBRiuDalilv8wb11f8htwd4I+0SbLg8Kv8ljNzvz
CItlbpqqz4iB37AoxHKFij4/OQ48z4gsWVlIlq4C42jjKwgQ00ESfS5cxVxUqSkoMRUnuPoK4mTT
KYRP3ngF6c5edZ/7q60ArDmLN+6hzsEZ/4L0uw1bndP2i/YJ3nNHSY3tM818xz+e7cAJCe/4Gtxt
YOM6uo9Rqu5c1R+IlXzPkZ6VHBqEpuKCz2mr6yOc49A7ybYMjQfUvAA006L+nSEbdhO44HZgozd/
uyK7xDqIUtcPzyLHvX1pmm0OIIfwyEwKJmWc7doYWpMmnGUPKfx4OS/e+0wq3ElklEIrdZYN2sw0
1jEAqwAcf+H++3PrD2X6jSSOaynruN1iJs0vABszrRcTYWLa1/U3XLlV17awXNqbMOtY3sQoqRNi
5j8MTRsKSZrAfHNZtG+F54qnIcCsfHhlUALaz7/5KYNtGtSxUlHhenAka1LkGL4lfHKhugP4fSok
WcYqbb6qADAAYzUscU5lOb+ehv2GHQdrIjt9n8BnuGsZQqzG08qOmS8TXvuyFJiVNtW40Isk5uY3
gKCSL7/VQ0B32uUVGnjb/MXKOrQ3kPsaWNnK6FFVeWlLE9W1FLeuBMEnWWGsbMiHr7Bqrztm36JY
q4L3Dvhe3QbsoEnRI1QZc946qMIFLIKfJ1pwyiJHT0r7IfyumNUpL3vB8vU/dJR2gYrvNgYMm/R5
1UiJaeVscbfswWq5dO39+dopFYVhQzFvjwvJp7gMEtRVMQTArnyzJUEUt6iTypLx+pk+ZYYANIjb
Ikm15iH/0gD7HxdCEXVNPNp6KknfGlgjLCtHj88zvPr5+qajXCFjptr641Y5QjeWrDUomHTVZMam
e7QvH6TxSIxE2BLnOgu7822x3TC+5t79CUoH6jQJr0w1gklVds33fKiHYCPLoBLXgctHhIJbSwN0
m7xkFMUKCFuk+hLVUdX9ahNbzz2+PKpdLYac7j6QBel4cSH6ZvjJccE3tVCKpv11enm94PTDuaPk
w9IEnGWukfXKg0MXMp2z8JnR7umRYEMiyI6+bvvMd4i4zb+R5NfizSI9BWdzqYTNqmK9O4ulaP91
0muIMYys2Hj3HpqHO9OgSZWacRM7KuWAKPo3zynOXGnhbRZb+RH5GrN6mABWhdpg+IivIICFtdAA
Zy9qK+d91SZCK8Z1rvqgVDFa1SEXTQkpiiKnvLYYJoPJ4p2no5taeiom25rIMcGn6CjXTG3dHqmc
kkiwa2MGRyu8usHSfGMs16BV4KihidB+MLt0cl0cx+dl0XGq6uKYbr73MzerqaXU3CgbMwU9RKm+
RLCuahZTcCBcLzHJVSRtTjG+1rFlwfvmvpnsblzwaD/6/Cf/EDSoGuLNb5MD+TUKqyqH2MR1qkuE
Q6hISBntzfiGs11im6pAWbsXk34wGDpqfsTbqkB4sawgxuS5LB3InY9BQNFeO/3KFSHkCOz390Sv
D4g1uLZ3aalT5mkEOX56iXrnl/ZkYAE7c0MavSADF2t4J/6sGNWgBPpV3J1e5U2g/N9D47ZYHPlX
9KETR/lY/86ch8P2wKnP0rQLrNKkvcmONxGrYEThK/SU8MU+q+iwfMRqqQZKg8Y51cIsHuoUSARq
Lu0r/oyK19SvMbWWaV+snz5/OptZ5hEW3LGqi4ycuJnQAPwWJNkeZ8AkhtRJ0WWWMfpwaT7EJmvl
/+ueRXnMQBCPncans3WI4TXgf0rnaFv55p99od3hPXgbao7rcZE8PMBhJOsFE4vZp+YL0IFZ5aJu
J/HbkMk8nN2PcytfS7ZkYgI65HTZ6FcaKsXBYQ4WQ9HMNv99Uu4JhbGKKj3M13fZJdQBfKkyk5a8
+w1d+4BUmScLz4N4XBs+yS4fkkqQprSs/BmUDeXu646wgNw61QPFiNA1xm1mmpyb62FUynYEDpn8
WyVw3abV+o3wGG3slWW1NrxIHXaQ5jcBWePn4yZSrouv8GaCCFdsEitLLDJIWqJflWebZDgPPaXQ
1G8h8gQGArSenZzkWs9XNm1npdyZkAGKtg47C+HqRmT2e7PrUA4EI8qOrd4mGKrhChny+TuXZrMM
fNGsiOb8HUcWitZPBXtty7+SkmIPZQBhwwvSwlCTya9vLTSRJpZCab+rgM8hZyZ8AY/prMAQ16Dk
L/Ekh1vVg7+5VHDO9yANcJcdif6Qy50xqXQb5XV+c8ls+6KWAlXVX2K4IL0SJHwHb60/RVnNNGwE
smvLNcSbFMWV/B7c/dtCruAkK29czUeVrAmTXnknSar+WKYMV0m+U/SwMEdoKoJPrrIeAJbP846x
abcX0BQLjJ6SbM4IjL8TQ/s/HyygwJQdGjAK0muWYsBDPO/3Dy9PY5qIAt1qNBmVGMxhXA2EELnC
GUT2VaLq/ol/R9B/j5IloORiScivxstgpqxsh1e7b0zAZzS6Xw/Njt0EWdGgTz7UURy+v6pt64J9
Cyx+FUF0rOQ5yeqkFFwpt9TR2O2QKRX73W9TSmt3xy7fngGgnoOfZOagWTKOcNN2B1+VohL2I3Nv
aBUAec9m7kDbI68AuzePOfPlFl99s2U6jdCVf48bArPd7y8GpmBn5bros/ZX3ENg6YrKONlPlTFC
YcPQy38jp9K2Pct5RnuEfAMIOjaUFlF7ZH4Xb4DWzik9RSb9FVP/i7f2iFphWIn/l4sPNkqzy663
hEIbQcmff4eBbk1m8aNC98PR3wqiwtl8HdB5oynnZ8kWvrueR8Ht+uMjWXbHtKlDsqjDuyICHeVD
8ke1sYaMEWpzHSKTL4TdMPaND5nYIR9briH0NpledoesiCr7S7u2keHjLD5wdPHK8pn3yAz5vIEg
sptD5HCeyLyleox+8ihEsdqBrt0pjTecTw5L4OMVkB8CfIg/p/GvJzkR5pbRm7UtbN6OESE/Itz4
V+tT4Xf5hQ6NRQXcgWOyxbnsYPPb85JMK4vEVh2AeLGulA4GpC3CaTR9xTc/qzzkMqXr3TSkr/CM
0pXpwYBTf7A4Mi2sUMjOVxFuppEvTZHnCKeUAsClpae4BEoqzE9IqCIKLYDxpxavWk1uZfpV6Kz+
Wf9lNIXo+tDoM5WEdmp6ZHsGsggvEVnj8env7VsoYCB/6+gWa7vIQHPjj4aYAjELflqlkT3treyO
3mHO+p+DAtT+lJ60L4smn0X9gN9M9c/RbPpTgELvRaPCuru2DiWLnj/2ls3APU9nq33cWaIWvBq2
qQydYFVexbccYRdSi9uGBUfqzetDWTx34U5f/mmWfBjJmK4j2WbMcwIlUrSKjhONlK8D2gZDf5qR
TsD9JvhUCPszyS4F3JgfI7sT6lBOKzncyzoOqz8/dLUycfIQOqe/TLzO0lhkOFV6wPD5BOksatmr
nzU0VOUeZ3li/4vKTV9y3cdLTfcJctjpMVDd5qUjCjwi1YgUpPN8QVV1NY8cLP+VGO21S/ij83VH
MN3W8Wx/OwkNW6JOsQI/o5cqLe5M543PcZUcwxm01OBLRQYe0xc7kP5Mec2fSMuDmA8bP2UT8DVA
Z2UbKhCFUlcIttqhPisgZnWHwcunWDfdX5P1ijknzk1FRgjGGg6LiOvD+shr/fl9znUuVTGaJo4U
KhupFjkr2LEEL1CRJ7Y8thFq8MWiUang7xVLWeeXOWn7cSW/CIwMor8Qqel3xDDukR+/EE+wLS/M
+KYEd9/qr0SStL8hodaLLZhoUv6BIHU3bZ3WVOVKj5Dexi/JXqAwWpnrnEVL6uwoiz+LPlGHQpC0
S8A6IdYIdZ91SMygk56mluvrnpxLEulWdvkHlzDTcv+GWQ6ARLbwj0mXXJfH75W16YvXZz6tG28K
m3PMYWZF7nvOWvt0OKZqrWTbTO4CQFGqqc+lEtLF32OSSafQhOEnEZCH5UXbrTUnzG82jaQ6DqvV
i/TCZK0YOnbD3NTmzGXMsl9DI6KW8+v08o999+DZMUCAeBKPc2YHC6IgVg6AvCt99CrL/+wZL7nL
9sS5bVxznA3KAUrS2AkNSR0wi9rDXxXuJX39M30YZ02OuYVyRU4+lcxdxCYUYxV2aqEHzhDS1Moq
sMXUL90IcbzPY7Q30m9v37eoKIJUePm4+nDOfuDPXMqnq8Yc8H+ubnlNAK0n8OZpdaJv30KDhL/v
qnDn6isVG5+e0I7CyPBjl9ZzJhPx5HZW7J0n1KnW212mJnuWp5wVyVQPHjwaPydEoOM3MbnSt9yy
UcmU4KLdVypgsg6iyGMEOL7UdrEoOzYGsDXSqzcPUgO77nJ2YzSNtBtCsPc7cfYykGJKDbiYQVPr
hOb3Kmp+nH3E0TkAWk6dGU99s4hn0KYvrFmmBzmOFM/FyQx+VuXreQGBSphoYj9Q1AAEmiqcpgko
rnY4voikkj0xbtDYTWr1o2QNVEHRKuohKcZCSAB90rySrDnXf2/fjASXy6XtqC2tDAe3pRCKjslZ
3XuZczSrDq+jbfCcPFXk+7fdCA9L2nFfH6u9PLia6ei4+sU2qN6QxfvOtm1ONtPTxFKAwEYsn59S
ky46pLokaDzh0jSGBu3gxtKchXPkKVXArm+cmucRmLPP9YrTFKPsKgGElMDcgBOOcC9z3Ph/RJ/l
4JZoOhJrDuqxVilVOcqPPopzZoXr8ReM108aZMRoAJBWyyfLJvZooEomEA0WtYLr/ZEYaBiUiF+o
o8INeCbEte8bNxu3tajKs2bqnaD5+XMkhboI+DEpcPjVfAuAPOF9DzkaRhwA3PUkYSxAu3JG8weW
Sw3IvgiGzmm5mRG8CTqTMW/zrUDJlHQt+5k+ayhdzOvGo3PlRBxho9dGwHKtZUw1JDya50yj9gP7
OldxB499c5QJg8/AKQ+duXW15sna2XoJGcpxwupa6hB6rXIxSxdEb+JA4o8g1epdQiyjgsKu3PxE
o7J2sQaWkezluAy7abSP/p1VrIjLLUN6RomFarVKbwu1O4mPl+UdHsZPQVl8ACCVnEPoHvQ0TCld
vPKcWYDQGw+6A9aaFH30NOnK7pLUhLH88Y6yAz44QBJLDVfnewebE6dfVOfH/hrmF03+BbbGBLIU
oF+LZV90Cqw8ZVpIsu5KDbvaTJ0aCtAAV5l2opgwZG4VqoXG/VBHzYwFK6nHxH6EvurJRiGj36s8
pqyjOFxj4+CQbqe0Jk3ebLVK1qu8bhj6+rAtyvLNc1NjN/demVZQwGyICATult4luu8vIpVTTWGG
eRzqsWgL0MLih8+SOL4CV69Gc4w6st0dogomLJzBakTfhZo67pY3/TEu9WF4nKZMs9poUJtI9PFc
AbomJaf3qb4vkqqCLlHKCu8Qch5d1MuEwa51HbdTeOQYSuUhNmrREWLm5v6oLYTnkkztNr5O6It7
YBX7mh+iATip3wGHw8h0vIBt/SIf3GR/btwvr/nNpMFwD+zLY1ulwpEAnudIIGBi7503P6LERgRG
XUjPAtytie+BBCdW9lvOXJvd33VvmMcfsyCXwMJhh/nHWemmKwOixYsryDu8S1cdNsezx+ZGH20f
2GqOMFK+Xu3klkMwZT8n/orc9rKEHWh9tiQwxAMYbJUJhgCX7RCdGKf6ICb5351l/a3Ii5cygbUQ
PqNKdPnQGh1DNAkJRtxhbXmS0U1RnbMXAJRqxz/CCoHYqX29Hk0ABIGBYMVkrh9PWay0GyVIVoWE
gk9MQ3FnkvXrW+Iq53codXtuT3AFBNEX9ZPfVBba3ThJpyszspYkNw/+Tjlr7+uaMKhx+lye/fS6
Td29OTrpBlGCK+hoZceGHwNYQyiG6BNl7/TaSG784VaUJpw8xfyPzw+lBcRPl7vNTnJmRRXK/lNk
0F0Gj5EsRcOB5C9A22Ahq6xa9Hf7n9PLqlvDz7tmmYlZPCnvPZLhdrAvKPhcnCBWYhNjWKaI9CCS
lh1aVn+IWnUEwvgdvIG2xYOSz9g5sp/MHVFtdymRWUxJzDm3+Q72+zXQbcSY7vaPAKm/Onx4fin1
Gm3bA9w8/WTyDDIWRIwtxqq01Xnz4maSsauqzK5GimyBSZKyfzM3AIUSG1Dl0lltefmNsvKT7jEC
xcLStnNmYAfGOZ2P7SUH9VDeS0gdb+4VTKG71JNrRuJUOUW/dERSdU/mewKxkCaqI8vJ7F+anZ4A
7LZNETg1SGbVhpPvPxDtppTpkj/iCcNwsRiSBhFdZw3BbUkPHEB/XEJ2lbIrfI4d2M+z0C4e4q1i
naHe1Wl1caPl/xFvVyLLKkXj7a76GOZ8Npbc0m6cwUpAtKcbPgPgNr/mMxpCNfaNPxHbRs2yLf0A
qpYsIPHbgsYH4sNOPDCHt1eRqO0SMr0g2mUIe5w/n2SeGWeUVjoUJN3dPL5UMJQPxC+tAWqk2y8I
EIhZX3IlPi+Fti93ANH11okMUperaPlcJFxYhfhDVy6yDpaxCoGqJTkDyUlKOKKEgbapEURG9HcZ
xfCxYsehvaq5mjf3tMRJOeTx3S/Pzc6RmNPvIgUDLYomHS8BRVODXHWRYWicN4M03+8zNA/VGny/
pPlhDHJrE4AxCEkN/oNagzzQCRp0eZQ1ujsOdLfhU3/xbMLy2034wA4SdpilWYULCX6Om4B2KAxX
stKC/t0yyrEeg683U6DPeIsp23oaRw9N3WRqNJ3L7WwXfHty9GHq5YcAx+9GenfL95z/HmOPmCeH
yOc6eGw+hGCexJ9/g8bw9cEZ+3665zzk+Fbbw+1w316rX7PplTIYKHXQ5bigbtHg4oT+faFkZK2P
mlsfIHSPQZTPoc1+Uv1Ve+8FU9UMr98FEtTClwjSuRWa/llBucTXHe7rZ4V147YAEwOwlecqafOI
UlQ7IvdOuER5Xi29x0Uvui7VUTf0HzroqKYeXQ8LBqJwH4PQruGz5AsWI2J8Ehw56K7mTZNIlpS3
lqCSlb5gzSu74zhFaFCQcomKh/xnrn3g68yEDRadQcpoZMh+n7xmsilnZJPJhLEq2pCJ1ErHhHh0
pmMgj7er9dg7hdkSs6QJp9R4L2AZIiwzgD0Qf3CgM1wU1bmai3l3PTc9+A1KBZgF8kZqXaIg+eCy
VikXAQSIzqDlEb+qDQKO3j8/1R6ut8dm9TRBR4423kXybBeLvT2mtokX6wSeIwadW/nxvS9HUagX
rDoG5yDrOV26bTHXTP9IrxZRpncH36sq1m4zDUyKmyFlX9tHPOQMEfZ0XnQE88qvDLhLmjtuIrOG
JbdrGQ1Sio0AU2iTcSNFR4Vv3d1bz/wzPbY8Jlhn6+leyqLDvo2qj6y0DxvPQhPluDLVy2uJOf3P
4vXWP6uhC3rB1RXCoYRJ2XSii4Ofkezu6GCqGiDl/AbNpzfBN3hz8pAsSaTMS3lk9pWQLl+TgjrR
joCu0ipteEqk4QAeVI/w2LI8NNC+T/MKsHMuUbymc8fB6Z3zxoWUoRNjfskQbgbXFtLzOL8HkaKY
28p2X6vGTTh0uHpM6Q7fKgMxTqwA8ncLvJ6n5pwVNtyEt2xtjlOA8ButyiNF0CiCagIe5HEW2B0n
9i53bUCPiSreOVCo/ztyJJuzZvKbQS1zahi60KBeuWXy0nfRYot0PTG3MLO8KDBS6l3bJQFwTBMc
xUxBhSlHpY7HPJziGUtK7FAIlQqMI4RSzWKkMnPypJbm9H2+b35AQi2j8zpw9PhWO3/m/f3SYMtf
zP6hghwURnSXvVzVMAJQGNSYt6mZNZ0smZ7GRm+G/ekyXESHsy/ZO+E2bqxwGZ0h4bRIi83o+EKB
zstcJKgtP0uLqX5IGnqSY/DRFAVLnK61qiBgWN1jPY5XEUtTOmdgWu9oIVWI50T1JvMC7EPFzOOL
ZL8gLqNLFWLbTMIWM9LIfb2nrTKbsiorPRZ8dw/L9qer/t7cWNcJBDplJ63/JQcMut2QSNZmXf71
PU9SVdMRZFP4W9ZuGCqQIGzU8Z0pLq2xGCKI/ruzkOTitK2NRB+bpo9rtvggQVrtSq/uvo1h2VUC
90LAJkds5VA/fwUZXli31PDEHa1iVXMD0fIQUuR+h5ydaPfp3iL7vazhF7OS5c9t79YMS51BYtAp
cKQRtjMxLD/T6obLj8bV/lmKbEqSdn+RQ4SnAJdoqKHSsxyu6QuCS4W/fikV10xfnYWFqJGdwWyc
slbgYMclbxKIaRNqzwdINRIwfL5HGBEPjqKNs6YxgfTJR+e03lpR9d5sVAP0nuTwUGAXXzz+aXb5
WI9VoQmIS+MdDnbawmrAZLssrzc+Eqh3N3u/2/cIZhLsigW8E0JQ7l/tcJbocmbhk/iXtQvzsAOv
//6kxk2Hw8/6JLZE+QM7NgfpFBuBQ2wNpf7EMkamEb59/Owx3Wto2ddkXMUipItFCV3fYNURvAHT
sNWPfnLzvsaS4vb75PHN7ThnBk44QSkA8yVIE5YteHs4ksxNlE2P05MSOKdz1fmfXiS+v2+g76XG
RXN8XQ3eVWhX26d0FIM3ybxdgzCWNlqBH9k5k5RHe87cuAedQyN5KfgfcFBqP3J9yW4hU5smiIUf
Od80ESdA9DLSmfpChg58L5UBcOGjlq10wNmgjhmt7oADB2mtVAgCjw/HGrJuOfK0Hn9LocEKJL7U
6r77S+QBzmRF1myV/DiL6rzH4vVh/qPYO3ow4Tnq8UZ0AdkLszUspL7bnrcv5TJChbVuFBpaNAwW
3Ee+rP8RR/gEFhSpXuFJQD4lot4UTJBN3xAmUNsQKDnfft4pOaG70iPDXGbHWiP2uz1/G1l0n64K
n14geB4QzEQErztXihbUSeI6JUtXN/xRDGLv3UvNVkt9DTvNjV/9BUzq96wxdtWCNwOXhLXO2fhF
bdQcL3TXZHs6DIY0qo8x8BOzH3JlQWP5cAKI0rez9ubZkQrKmhKleiCxe5wm67XMfe16NTsPX2il
tbc8354o8kC/KHyWFAHjZ2bevXSw1cseblgKqcBR8lpGOOySVRol3gvLSiDWe1HHj2wWlBseQ+nO
BaCQpaLx5dld/+Ygv9HsxH+s+NzrKA3tk4tAH0Bb7nkh9ljuYKz1zIxBA5F3Nk7JFUxLRuuALY4j
VvlW0DuK3fAkcFY6WssCEAIDxudSwYsMGEu6PFuHWmLfaCKIeQPCz7dZ6KaEl8/xvLAq84murHUZ
sOD8Qczuw8tq0VKctxiGB1SxGaWO2h8Uxd6pzH+BnnttcXnTXP9IEvHoQ1Z6m3Uuc7WNb1ksEL4U
kS/PuwtFIxSGAM38Pg6QQTJDOfo0eoXn38nXqheg1CZXhnEjbY0dTQ3EJr28RcVodzUS6Ko6H1Ms
iVCIQ5czvan9KGgAQYvduuW7HVQOhMOWBlIYyh6Ml7Gy9Q3rcwqbiD/OSFwimMVdHc5kHXctm1SH
snlcd4g5y1Dgog6rBqFzONQ8Sn2tmfiLzg9ioHyDS000Zq1odQHVqQ9PQSrHw/vxmZgVEhLPD9eY
2khRewraCda62Lmq+/W/KS+1whoDX/Bt4QPRpHkjepuG4Js0uJ8wNRHoiO+PMWNbb9+JFru/W5T+
TnPZHmzOvsNZQypzIzN2TyvI7W7Urwr0LzifL/Jl/qXQTRXglS0aneXk26HtJB5Ha+UHNlPYVIk2
lLU6hQvPBoV+GALsSe3TOTHjfMsvRJt++n6fwFOwhJt+QXjVXcR/RDfu4VOP2ntDZykR+54nxyWU
Mh73fCo7NhoDl7t1Q5rnoOWbkbm8QDaTIfpmbDqPKiZYocLcjnkt4F2BOR/Rg0SClOJNTYzE+mcv
uKsa8cezM/h7yJMKKYRJGnugHGiS02ah+/ItBKcnxgxlgWbAIFhFFH9GZEFh+GN3k3LUKM3gCDIm
ib8GJ7f4gdUYEwI75ULqskpgOJKbP2NN2vze7vK2xBhmE4gQGezIvMxq4PqM4k6m5xDzrLW9lmdi
6YSn6vD0iEr2Kfw+HSQLDz1hC336QN/TROJ7EMVPLBIncO+ZEK7MC5eXLsBgi/vFVJrIZGMm4vE6
KyPnZoayRo+M1EF94KaKCPt5NswobhWvNGcjKdZBGhEPCQ/Uzrtu8apvdvGxX+OCFJ3KxHDEXU7w
LjQYcOxIPc2WhAyvuNcKbWgFDV/cVvbIi5QnCSjn93XMXM5aya0pJUjnfGVxHhVQ2IcnggIFAy6Q
/ZQ9ja0CxDsSVs0CzX2F+YjDwbyP7qS8Qvo51VfqzG4mTBVf0qKHXVWg7v88CHseWiv4WGZUvUXb
2Q4B59IXBD9ygIxo42ZGKAbrS2ict/HmDPVoxx3Ybk2+V0kkj4nTsszZThI6Fe2w76u0acRt7FY/
zl/cZrJKXUd4zZDWt+WBY+CXlBvjtitVT9o9t+ebe3Kxz8pNusEi0BMnzvwoOUgXn8+suTwQTLN8
FjGS5kOFDAJdg3KOnFz0XH+4qlubusCQF4eWfLEVs5n8bXE8HGUX3zPkSAblK5MqMx7id2AMW75a
Mfh2PfLA+JwEjyZ3BWlJ7yBKD3CAM6tvh9btK3EMFLnaZl68xX9bIJOtoFuZr/3jYKgimOAC58TI
f/cGYzPSfGdJ+xRWrqLRZSEnyofvPl0JucIiOlEynk6LHvhIYLac9TlM2gRqnCKiDJQqtfoF0Bj8
qfpyuXU4amFKzqAZ1mgfjs35d4VQRHSH1mTa0yDnYo71U+6GyV76G3mRpru3hvsXLhjw8JFm586B
0JwFDZOpGAEFKMPOs4SzDBxODgVcYn/i0dw1oZ1SYIvHQ5podTYb7f48iNViy6YMJ0pWEH59up0p
My6xH/iQxWN7Ar7BzJJB0rZ0Q/NII7d1vyFFAJZbzPQXE1xwb++/47eQPDf+IPzO8D7LLMdak5IE
T0r57iBv5RsJWl71JoUh6o5woVA5HCq0MQGJKiTTyxgRdn0oR5AB5QJPAmfP7oaBEqOO3bWH+Mo7
88vOwXO8wtYFXwUc7Wdmy5Gwjxzy27JyVyaw4szq0SdDVCpTYw5fBc11opfF6fB6uQIl84oEZ1EE
EqLA2qPEWC2WsiLoBqSRAoL04FKIQPIExBA8azjinUzEIrxmizrOWHQDhAU/PLqQsRa+sq1d+ox9
KDOC4CY3ogTlFteXJUVgOfVdkKQ7ZRSLhLzcSVWmllmafnJDBB8RRnUFfM7itg+2nHCKh617wvQH
N61+a/0l9P3Kw9KnjwGDajuNi7a7DmoNSbgec3o/+7V783lLSFwR1OeQ5LCwYXiL/eMsKiiA/t8Z
y2tHp62/rB6LaHwb3XSJhFEhrKXjzst8IGbSC/xS41YoCbW57CMFj0sM9dMgLA8DhdTGEeCzycXo
K0qQUTSSnk/ox14cz+xfnnZ/9bZpkOhls/kEFHkFlZuD+zxlDaCXEyrvpdXGaHXh9uaYq+IYdK9N
iYDJn3hHR6HL9dCClTjmoV38hJbp9sh94bn5lMP8NOAIohrppGoW22R/DsS7oKEysztC2UTW8hMg
rgJUF4Qqy2m/j+bQ6OrEa1fiBpJfck3aKBpjILB7oQvr6CsVp+xQQWtrUyvD9wdaCfEAyvto2U1E
uyKF6G2RcYXF091AtzjKekNj2clFnYEwc7kcerOq8CZKdSZLd1AYWTKDbXBpEjcA2DKtc1fcvm5t
I1254kK3UlkP0LBa3k9Hs2qD3b5SlHYlECXhnGlJOtMLH7H+arc8x7REUK4Fc6cDN5NXvKtCOAyn
UleUR+UwVO3QwO/HnPB2cfzcVnmaHmlATkTCM2jxLyb/1pvD0EbRoWfB9bRgE2dz5sbhZdX500vr
StDAJ9WhIArO8Zpe6Cww4bxDK+cU9CJ5uePnppJ/kkJyrixP7WQFZBI9EXzhjifSFsSW1JL9FnkU
/pXYQ8GAlP1KDLFjjbrMY7c9DuT6/ZTIXjB0g4m4F5n/A3fi1SHVe52BUn6nIczOjZ3/OiaL04ld
fYSyGVbDkmgg/HsdUcxf13fBWUNZ/GVtO00WN/X4qgBjsDYuIcJzucHXnFo5pczUUWLKOxut2gEx
0oOqytRTV6+RtoG8etyFrf2WOmiQ5nRfKxUzKciqHJnki5CtOVCzWcMoxUreD05ExejFLCb448RY
EY0YnH33UEl6U1RSsJWmRylg+TZRcmGS9y+xxFkT/CxPTd5ki1tGY/4ZyJ+Dobiw8SORuNQqvBND
GqGC9VFqfsJ1NmQiVIX5t968WDPthUJQhnBLEXg0QT2AsFVjYUm5BsaOYvuVvQqC6ELRWa7HYP79
1nGUtWPYfpugCoED1HeFLDh6Y6WNzv+FqY/tgYnRaTVS4GtAdnRZov+gNTzf1ak2abe0vYmQ/LCt
3Absw/+f2p00+kqXnkctWAeFbxtc4hoz6Z37X5FZBJzfLVSBEcQkriyyYst9HdPniQnQn+6Ni2+m
EBoLzZaEhbg/fKVrF2s4WoCyfOoTqI9Vr56U4WpDnQm4nWRjQ54kpTchKwxq95uCIes2Fz8xlfXo
stq20viT0tzJPKghYDcN4Yi1N8AOFhBHehg10ZPNzSzgFfs02d8NUhLw8LhmvByjtl28qHbW26D0
Ly7DmXskdDqN9In/XWnK/uEGFL3l3JMUPnkreAIX02yMBn9kW7JmPP0Qk5MogPP/PuIE0ylH+1dY
0tHnZ6WmaCAb5bcFDvy1XWtaD5t3CwdU8BJxW4zzb34V+pEGPdR2fmoGT34WWVl8//u3EUiOtJhS
q9WATphXx9Ulv8P3uuTeC/Thg5AXVR3AbUO/J0i+k87n03eDdUVDpPKuBF3FddQblDB1cSHV40Te
hz5IY693Us8GLb4vK0LHZ6vAENk++nb0Qpp8qGW91SXjwS1eT0co0iRZKo3ovW/afTpS5Z+i6iaL
Tqk1qyqp8BwLX3j408/Ba41AmRVy51UCyaKH582Md/2P/rIUEjbFFov4aGsXSrYXAcqYPNAAEK/l
z+oxha6HhN/p9/idkGaRGurhKoY/iXhVbKRHklYZ5YIrqa91b46q8fyLPOB2WUp9k091A8uHpcjk
8SjZ88gzCD82msFoGDoS7ioSO9SG/H27oj94rD2OvxAVe0jeV0j6NsHeEA1i13TPsA7TX4IdfBOm
G/UxpZjDxSeUPsoDkkqsRejWWSarknoPm6mMw3ImVxXK6+wDssntHFw7tEKMwUGWrCV8CNockA+8
Y0d0rYrzdlPW+dhELfOnGsxOqJ6oyPXADa2/tzTMe+9HsX+B0waHjW7mP037HX08W3jX3AJA1VAI
V9Ikr+LxMkUo+bdAdhjX+66hdwvA+LZpGqkWxACkblpwqMUZYGXqO9TPmX/L478w0C04gS6Glkgh
3P2Q0dL/hyqYSLrFZltOCyGuibSt4oC1BeBeDpLSP9wxK2yLmxtlMxnYLtwUin/TGHkXC+G0TVH4
kC8AOIhVnegIqthebj4fHrM8XhNA9Tebe6PDlHLs7cYReZe/EQBHHdLwKCL+750ul6mRvAKZUErD
DdGXKcLCEcbBZz0h5jgzuZ5MKtBPPFNICAeMgeb++jXP6x2QKk5WYo+m4xjjCLmct1e015aNSd4n
GL2Yr+e0PN2s/NmfMhO4nDDOH1iv5611tH+8mGm9rCF/nyy4Ppk2YjujDekNpgya6s9INwnBFKn7
jx4DNbrKy4jij7E+03uQ/2TSHGuwqTT+p7UrbclXbpu4GFxzD4ri+KHYVMSrD8mJ10Kee+ybpG+/
jG2bH46nzORNIvkMySPC3SUTps6IFCwZi0K0rQOVFxAbcfYI5xgmJe+u7FUpDTSiJKqrOwclGsJY
7O3QutBsKtU5fubVNkSfSe3oPO9Sa8Vl5LTGlg+E60IaUevNICNMBJLMHA5U+zS7NdqsRQDqyvZE
ydmZipf7BsIV2a4fkwXW33FQ+PJmeJHdm8oPhCTMVCK/SSE5n0IgTJnAaUd3Vs5lRKicMExg2AkI
HU2LcVJIdD5TYpe00tdYRdPO8L5f2I1KvhjkXQmvVcjeYlzWQD2e9+4pab7HyzHX/NsWE1pr6i3i
HhDcM9f3NgD0P4DlzdegnrKGinuuTxlw8wmhkCBoDg0xTq+fGKB8VAjlCJQ5q7oBsxfLcv+AcVBD
NxnVvY3iFSqHezj72sXO/0lX/brc7I+Ow7hGGrXPEaC5FZFxenql8EfSCi5cWGINRiS45kMRgKdB
Jq0Z8ftsLPI9H2l9qFoO/2j5q8a7CiIUxl0XRQ+mRehoSMf5ULWX2lt51S+xTqI15qLtF/3acO6w
LzWHrLO+GabNgQLjRDCUibYJTweV/5QtezIpdefRqASaNeOhWVDU3wyW7EtElyFhUwQWl6Lc0TJW
TqG0xHqVvklNgG1eMuKh5CuD57gUy0HPb2hJwnL0PPZNpGzRPueUpgyrDqd7nHJC+xEn1lWkrGly
zIi40zhFbdRxQorqob7EAsLGlHicWW2fKKrztd6pyvf4N3C/jLQJRs0zishemWi+wWQolFqqxuzW
g+oSpfY7tlefG/sYrbILpAHYuvi5wQfB8COfa08byrTu6wNd7N4QgGJZ7vekiegfoei69Oy4rTDW
MH0ECGGUsWjAUdsTGyhvr/zkd7lN+AhNNQhtre1O2JtDZUUTY0843Pycpf9y2ommw/arFIaQBeSd
h7XNjjut2a776Pgk1+wIqyR9AcxOw7+Cva9udARZh9rhqr/k5K2+xu0WaIQ9zyyBWzXaRqkF1OMI
P8r4Llr8m4TxClB+nhS5m9UrUgiggmcIzQPm9oiLZfCbaMa/N9j3lgGdqCJSOPnOT/3rcJGTzX7A
WUUHTTlXBBGkXPTMOwFHiofTCufB5PepUHlUGT2TmR5t/TPmlFIzjP7c4CHQU9mM8BS1wp3qkgCr
IUA6zBVdrJNlxcDRusZzMpsj/QOnnQ9I66aiVRGvH7XlJlSrhQequcrTVefVNzxDTI12JLtQF/7C
HAiD1NpTLUGMvDQr99f9TH09zoYLXd0BLQu7yQqX/KnMcgrgLpq8PeN3YQZXGZZA9+ySXiWhK6l6
RgZJjl70BbcQyjKZRaazaefaFR6gNeQQV4gMavZI3mOIpxF5uLrodqzU+HXAKPFftjUekfBBEtd0
tdD5Wz04QNv88IY14zlq+k0RuV+KKo/VaT7ztuEWSVm1c6CvHCQXKpHAVwuFT9vsN8qPMb7U09JQ
DiaxvDycQLTtSYoUqo0ehJ4Q2GFtRg9oUPUl8CH5oL3VAedbLXBt/ew7IDH/aw20s+9tNcdGHl+x
D9OLnFbdSAjKKBA65UnxXm5yfVbxyct4YbCyyj6JTfG3vWAsVPiaRFkOpeF8389brpwD5HVtXRZ1
NIinpdU3fsXFd9zjEIe6rTgGHrPjMnPbQWmba9Hy7gkzLFQuSHSNYZF10WD2bu2H5u3uvs7LmQr9
PieSiKs8sPwK/t/MHDxzzWSgPH8+gEiuthwlmaRGnx1d1Dnop50uHjlXuxYBPXxmWNBBWQYD2Zcn
nI5Q6JydlmRCgflWZuvFJaqkl47h8EZQcDDOOVuwkF4cUKsgCAAHuEOOLDY3d2bT8egaeBCvkxnG
xOMAE14P4XXXFatPYW7oigodESEyImUPeFB2FdiUDYdjyslo1g6krYvqrAKCkTeaqdP8ZPc3OZ94
ASw3Q8FacsEfgCDmwCifxxJrTDj+Vq+FuOVypR+eaTbp3JXtLndl4gtOfFW5jzgr8fTDD0p0cWz4
KwBGCC0dBXi/aJgek34B7FUuhdcqSp2J13x88DAMiGetFAKqr+ullaeJ7OEX3fUTy253V7qryK9Z
KnK5putPV2Hll56rNpjT7cgoof27JZETota8/Gwz8TvHJAIKnObW0udyHVVpF1y3PptgEjppNefc
H71Jt0ZqWv7Ku++7vS4pawK3xvqqfphXMIcGTTNtwB9NHUmDpQ11KGLtX0R4E5Ui9f/8Zb+YHLZs
rHuSGELSXjDIzsHNPNrH9kB5HfFYWiGS1piUG4jCofBrSUZl8hMwYis9qpBuYJO3QT19AT49gunq
WR3eggRls+jhDvM1tk8U5H6Yy13eUAvpBqX7XsjMk/HWW2qqJTmsawC6w1F3lpdi4OX1UBZgawCD
qcu6l/A8VhRAyBBwvbSVtwUDDlVn3mKX+4aZijSL1hYjmX54uMk9FXlNUuT496o2bq2Wzj0mLXEG
tzrjq6ewAtfZSkz+bRQWGdA1C5v5eCUMPe7PQS/rXcllYx2yl91ldvl80JvTNGC6XkI4KUtvtfmj
/ss4qMALOQd+98RQ3ppIfdL9l5+NvxKVhxzdpTQ028tQ9XFLeR7mhuFx5XP2bxukb4DZ4cRglKJS
uqYggjKlvVV6xtnmejaUlkhwmD54E7cUNWCnwrU6qkHWUW25iaVCXhjeNV4A6gmsd9ILMFY5EY8X
zWnb6sYdeG4YqJemnkkxasFtdfQnS8ixih+O+OHqTwnYHzG/xoknwStgLS7M+3Pdy78c4p2f1UER
ioncISObJLvH+D6WMAdyxsB3uboA+QEnExZ10nYnDLfHa+TcZYX+9KLVQAX6RewcdZ2+xXaJE/W2
XrtroLW4x187RYiTrIOSNIO/A7pYm7AW2AAdzEvWaR2ZR+7Ax9TVDxn1RZwpRMxApvYHVm7AkuNI
7L+NbyXvCX2ONop2I57FajJS/mt3U8wvVCsElG4ywsBIziBGpN30DSHB2ZZvJmr5PziMUNxHZZd/
ZCgwfxME38hVKsp+SAbldbq3EqVr1M8tGY252ASCyHCfln2py8SdIrdD9SvJys/plQyl8iaU+TwU
jTUHGbInHgQnA34lMIrCxEPqCwK/QLvkUIv4iuDxFb0s/yl14bR1aAV0ofHe5tjCaUloX9CiRh6+
hrPWXZBtQ7YyMnVbYzcliW6hPtS0DEb1g5VGLgaRWKAb+8Y/bTVvMITgDaE6Lg2Ol9DaNiJrH4jW
zYgqH7Ewg7yzKkjw3V6aO0TqMbgw6M4LDA+6JmPyaW/0yl9de1d8iLZoYa7OLsBc/cW9KKbcpvkG
k/vWEV+VvgIStliL4pcOdpEgDJ+iEFdYHFUpAeQQBs3JtlSrO5d80LuwnQTKAbE4oEP2vBCtUEB6
iNIG3Onas0660S60zBtieEwJzCP8xA5sVkbV/Tqh1Mc2Jd+XHtHSV+Zh8uhKgyaO5Jz+o/lsMZmn
6bwrJYMKKTJpEBy97VwJVr3SPOqHWCParObQzR5Nrhne8OLgVGlfOU0eMdqprIZsTh9ahJ/CHOIw
+YjK3HPIoK/uedm5aGEWQEriS35d0uXqRIiYPe0Ti5Ko9f3GQAa9Fc9KfrBe+XCmU3mQncvL+S5b
YXGv+QGZK+Bb/osxyABh+p7IhQKH1lFrgojgjmuREcemWP0RGpMsOWpx4MHDzt0r1UfKgovpbuOA
0dL/NtlmzoZ7mc6SEmdRLrFWhq9ftDBMtWFVanVCxQYAfU4ZO03NY26bQP08i41NuLvwIt3jcbk7
zpzl6IQP3cRPQRj4noDgyAu/V50dvArsgP0ghWWN8I1pDllAYUNZvFhSWFPStoFAUnjcmWze9Niv
jacrPYJFPo2QMUymoWMKqwHZAHSo+c1ITyGpkEOQr7kTx1nWiiSw0IqiRO7AMbpb06Kj11iw08mn
PwhyrOtrLeHcxFfRe79x0nWnW1RBibGVBzudoC0ZIIKBidJ4+lHBd+D0u6pXg72DIFsdqUlE5A0+
0m00/61f8jSjH4saVKLOLQ3CpM5w8n05JBTbp1bsi00xvfyDa+HuhdVgDRJ55pgkcOcBhIKjPlkk
UvQ6d8AZptg1KIPFnJwx+i2VpumSDvuPyRvRBHP8H7jMIURg6N/gGOhpJSIVpx1OMUxotqalWs1v
K1G8TacVTw5tnQ0LEn8wobFZ50fpOTsdB75xmmvvDhmnpb66pFbf9mfqGFUoOwtqCt2oF3wQhyIm
Yyd7or6rSU/NLUSAUGFlmu0arL+w/uk1Hy0GVx5z9CFvi17I8OzLe0ioqxSfj+g9svWY1N7DbwMO
Gfh1E9GwweeEdhYSCUIj5qH+hAvgJOrTmKKkOsESLj7C+ZFZ4XyOhcFvwT9pqtN8KBVlXPIc5IOv
6uWYG4BOipCkevnav7jXZ1WGbRufeBEaveJiU9bZwLm6/6WN0acI3xksp9SY4Mt3CJEJoQ3NLCN3
+CFx8KmKjeMGzPgyMdGRv2B1+CalrE8/2Mfcm00VuzsLK1CHW+Afy3lpGBxr2k9pDR4hTNsZPsWx
GDg5aHC3cI9S7us5gUCV1D9DK9k9o9VyD8M/qzX4Tpk6yyUXkedF1KcqSN1EjfFcgUvAWZZggp6G
B90cTgwLTgB/3GF+G8ec+mvHJNTJu02VUGgxq1pHFyY1Z6QpsIWlJCNP05iAJX/vs8r8HI3fATM4
Dn6qVJ5eFlIQxP1S2yXrSLeuPhK4wjQMxcIt1mo4rEYt8kmsY5eOgNaa3gqO/+THcSUCWnBxAijQ
naQq2WCT4vgsI70hv3SteIMCi12FAr+w7ZD/LTbJuzRjjsi6H5Vyyw/1XvOb6UfGI8COBdp12KY0
Bz8IUj2hFb04Pss1MF9hUUkbB70e2uzWioWyDQstHoBrVw2U2lW2O/VnorqCGiSQ5fxZ3L+2g4d9
VwMPTGhYeGSOFGFGV+coGjzKcrAuzLfP5cBUZziLBWHUtmE9fMDk8gG1ZtCf7aEkgfgf2VCTzcSl
Efil4Ol7sKJzw64dOb6T+JaIFY7Y7lDSLUSUZzJ4qxd3bwedaHETnXFy2Qa+TrrSI+9CBn0ee8OM
UERZhxZNEvUaZmIdpVyOlL8SNOnihCoY0WOHGzvNB6heu0K7P6ojA1Bclnxn3Jy/e569fZSSM+dJ
RSobmaJwtyI7vVs8oW+I/lGicdyzapXEAUn+6xYU7Y+6xBd20YJrCOiTke3Dk0AMbikCvvxljxp+
ZJcdtAl3EZbQogxoZaSooIHIQhFg+OhoOfKTdevKFNaPtOY7zIDtcdO2jJPfE3pkzH7OwUDJw2zd
JZb4N00u5169i0oVhMbercnLDtTrDXFubrFXLEazApxdHuU/evIYo80TKOv6qeXqWq7Zhor1WfXj
GN0p5ugNzto/7ZfozsIFiXfxzXwQQ0mIPtE6HIJ2ndJb5CQhsAn/LyBJYu3bMEifTLsGOAVnCwmH
zeCfox89NUUlBE+CJZiwLEgWNPf8HTLSGTHGavFk9wJ2lpZ7Gm9N7wPGAs6UPS6HXSML6LDBiIwm
hjm+bwpwQmlQAn9azrilpkUwgwYLCWrbgAtnJqcKT/z9Ddliuym0FoWLkTAc5goU0H/1H2OFbqaJ
MG3k29OK4z0UHuUWZLG9/6/7LTjNn9TrAhPaAeaGK/RAHY+JPpkwFtmYizM4S33fa66yRqJaK1bm
ylWhVoI07ga1OcYuhyBiiAv5EnezvMSso9ubdd0skQt3F3UUWOyU4gSx4i1XMlmxxbTKgFkLCfzq
Hn6KZCk3E6zbVDtExz8+4It79Rc5InuPWNVXmCRHC2ygwxp1pm/6jUlh5b3m07jxYbKkhWPCwY40
gdorxSCjh3TwcSTOZXROnClmmFPCQPbY9/rWS260Zm6I+stv/2woAyyr2qA4TxnNebzyYnw02cx+
r/zeEp2hHKxY72Hyuq2LqcfpduCUwDJ2UtHIbI2gLxQdBl4z6iIuyHXml/E1tT4LzvCaOCmf1pZZ
G/jWuz/xvqM9mXPAMSbLFiICY0gCjiQhbuPkkU7s+ysqOLozKX5l41SD7eUYuXGCaLjB1fVOy4Na
oF5FYQuLIMgDpgRb2JV98LYPIEn1QGh+m4pWRGRLjnGCSmGrgDShwBzb2ytwNNICHGbCsIDmoAng
qh8X6axlhiNCj36Brq0V5RteUyJXRWKIgE/mamG3N7CxdUcnfc1bQM2oOQkR7gJ/qg3RU7G05GY2
BFPc9iUa17HoFh4NRVHSC0EAwOAt0Ayz0bqDxpi7EBhXPv5FRMzGSTTuObfZvpewFAEYK8flMiP4
wlW60o5qn7p+2R5s82iQZB4SUH2sLJ3JU2X/9w/GJrjKPBtUlYYjhk0aj3upnYOwu7ZH5KcRu2Nv
FTIX3+ea9nrj+6AMmEvQWHAcxpaQbpGNzhliGmVWoLZOXVZczYJFFBCA+bdM8HPaPYJ+ylsYC5YU
McvQJsCPG59qO4yImN27uh6+XPAfx/TuAkHoA3J0+isFaDW0jU2wYN3G1bBnpSNA6o32drwwbxKX
nuUTFQx4GwuP0F5PvvXyXH4mSw5HmXA439fkN5z+J+kYPshZbeHEkTqCZHAf13nXf+NMhmANWdpu
C9UHrf6TupiWnSCJC1mTwEeZdbMPl5jqCa/D1Z9+g+C74yjcuSkMFD1cRgSYWtjzJKMNYFRq/SBj
FX3Xr3Zpx3cwapKdLx6FMho/6pE48F6LoKjy4pODZz+9Z9ALelVmkRkJ0tnaWZEn/NGccE/Wwizi
IZE5uR6yX+W90NyYpiOhohNhNKPtzpgtYkAwGqk+gwTfX1D8A+WKhpY3yMawGyeoCRPOrRJ5Advi
bC2l+2nWx5mBwX3rS2IAp+GgaTXt1jy+aV5VIVVYym0nMFcGSGhRp92Q1/XxgJGYoApRGJS7mfA8
KabnwKtZf0GZLf1l4Lls1XpB+NOPS0+Cjf6+qBOWuzwnqJZ57hg6uoQSKwWPd3dEm8xygqKVOpm2
FJsrM0Fzq6K9XK1wsNkq71AiBXpWOMMTlMeX5PkESaDEHr7JatzUA66behjhIGcL2rfRPkTzR+78
YLiSIGtWim2CXHimTBEo24QpNCuxMk+Iqui1NcC71b6K/klyCEYhK+ahUxfAA8MnAcENqToWeyHv
3gpLdH0IwjipdQylloYvqXMSxMVuKhzx8K3AgKrRoT9p1sHde4xv4JpIP/dkLQcYP1iphoxRaOS6
ENdzMZN0HCIxalWGz6mQNMCUSQXi26crOzFXwONFNmBuisvyTBLavbIOPgASqIt71UhjpyNonc4M
GtqglS3oT1iVuufQ8jTpI5oUFpmKo+QklyhJz1O/v8Xt/aydF1PvoNuYDsHlp+H3LaL0ApiobhKD
CaNcA+VVV8w18ZxICAcCltcFgSVuG+8GksqXp5aEdPm97rv1M99VV+JUDvmS1xJ+LehgfTfCQb5S
lT83EnvIOZgPNp7EyWdy+aGiTttDwT1o64/8UCpf0mTyLpWLfOVAnZvGTcJlM9DIlblVOdpO2qBl
89zYWS/Lm2De5uT7T+4z1iAL80V/up1Tqzz111dJqDW0VeAZv7jk/zKBls2Vkd+JulK8ccpJ81qM
+yrJ2romKhKYrVZj/Skkd3WEDrsjGdkA4DWbtF4n0t35AalZQXsBfZNw2RKNrDcamkUwLnjFwfSK
vqGyxFfQzKruwsrHsH3UZ2j751wdkiwpXy4VZ28CPLUVJ2kGPIEsq+OokdxWTgv/3dOGWMJpU6Bi
J2h0xtn+Qx11qWEFfXuzRdbwMpfdRFtGVi3CLiOPVMtUQj+Htqy1gVPPOm1AnYfm2QttXhI38ZtX
dW/p61dKbH1HpluxiArjp4LoGZlxwPQkDG8+VfFKY7/9HMS4+sMZDRaus/AKSLH9PhqW+6hOQ+pO
hao/+cybBFa69OiF8/pBBefgAA5UbdFUbKjD2laL4gTMrFE5CgT04KeLpLc2qIKi7JH8QDpxggyJ
RRcyZMn72o85MkTxxLc1zkal9gfGQUGSuNaCtjjSuSngId2ywJ3LM/rpvxZ7rIYGqDKqefjiwlhq
13SVoh+UAL3uY/YJkZp6UOinbIqoCZafwavnTqfMoK5wzf4395XEjLOghceMI2C6dO9I414EQjtK
uz3BZvvRG/KZ8wXJpabUjbKNqBB5QvUkOqxQCZhlDeq/9AYC856V2bl8hu0aAdDGxIINCybpnEYr
MsV+HRnndB0JJl3JkYAYhNgGpIvOJQpG16MmPXA2QZPRwzF42TpcENKPV0al1GGA51y92xTazCkT
rdSJOCWZiod6RPIOnKzkUtbi2YuVXzYlvUnewv9I+eX2XREcF64Hy8PYwdp0q/yDvaks+ZcLfgNi
yVBDnFQK3pnNxinMN99M6LbRlIMfV6KefnoJsPcfAyPcWXvxydu/KyLH7E6XtBqb7TkhSNVLDOIe
4UsdOyUJN87TVft4SSHKArHgjKMG3vCLdt3HJ/xo841MW+1vmy7YPYgiIqO83mn0GF/ERgodt903
NyoUjmD4IehXYs7vNhFemfFVNxe37HpV67f/nvU+/Jjfx/HXpHnRqo6hvaw8E8pHIQG8z35ikBip
kNhV+TZtXdu0o5bXDwuLSqSJgg9oohHdmwKn8IxwT67ofcQaOl8kJIuu5NdbWviSkrVFNbLKkzqW
1mQ3HpfeCorGxuSa7oB/u5Fad0sjtNvXcUMKYqanEKR1mM1f3ej0yRCNn1q0sujFhIy9skofnFv0
5RGnGbe7NnjbdEdLG0u6XuGNpmI5YxDWXtrI856E0trE3HcFdVjbHCt+uKkGSn4f7TCCk/OJE0ep
z9MfO9vuILT3ZBLB+vmLVOMgdC3YqwZ2X80fiM6QTbklKCJ9lCDju8B47gdEpPTrM4OQN6ts8smN
VBIgoQ8lo8JljaDRjOS1AHYDOw/y+wf/piY5/h0OVlTfYTNH6JqoxRjgssvWWmFrJoYiMSOi7HNL
re1TZ4KQYlDH+TGvSGHJUPvgTtN9k/M5xasxWBffzQfwcVFWPOo6GwLbXEKLrGZVQV79Dipyb7f8
t2Job9eFa+CyVgn4qGYI7Q3Mfw0glc/DhPFiC0gHcqzC86fQ6sPMNz7VQBTZzemYvApD3EyTGeG4
+S5rdnweKr6wWUsdj2PVPNcF1dAPaOOCROir80Cih+6p+C/lldyE/LggyzJG0zNByEX8mlkA2jWR
RnG1UOs9GLAVRXQcQvQ22zKkGC5vuxWEkhCc4kf6YNmaWaVdPKYrKo5Atn6W2lH2w/iII5/r5GZi
5olJSfk6/TqKcpBpf3H9Zye5D9kn64Do007W08d5mjGvwhF8LqC2LJ5yZsf2rXixYvZrvEG6psSZ
QIiZBY9wVV7i+c3yUlMpSR/3lRFhxSG8dD0JoN3mZoIX13lIwFY43Z/LhM6RtBI+EraI5bzBfj2P
oy2ezOYRyhQfVg3XYRnR35qI0g2DxJiF/5mZ105Uu9TGIGd4RCROqs84lydVCaLwdnEh1hGmLOpO
ysE9lckOJ05wCfmkggSAYMZySsRqzqg5hUkJqhyiQUiSofzJOdK54AYG1VMSqTanxlU/GtE2OId/
OzFLLYXyssA/rGV0SdbZ3bU4Lav9o9Dkd3XREKtQ9qHULHnoFSfs57h9OxZoayLTVDnzDjhXlPAw
dQt1KIRXLjLgX9voyhg1E024LWX33FY2eZqqnFqIHYcxjLeZOy0vbvwuUXOvLXeKgwPA9BVwRpJL
MxyEPzx7YgvpHvYsAlXbs8r1fyVcfBaoz0rh86vGGVHpqhgv/AgoYeHKQJ93EP8UWcFiJ0br7SwP
YCcgdSUGlrDHzZ2IXSBF/AcWVAEGUwHgeXl7R9qeVLTC9AsUrSS6uRpJMI3B+4zXQ83JubpszxXH
r6OhRO0ydY7sgFwB1hHlAQEXZxlZ18vb0j6AoXWR6GP6NMKtjUVhd36sQLeyG6We6rktTnpSb5FF
pAoOqBIYctsKWdBQtdcx4VeHsonMrFEhdZWS5UAhIMv2+k9f3lw7z1vQ8dsuOX8L2E1QaGYb22Do
gtT8cuaTjLMJQB9/7b0+avGNt0bqoOqKUJP5asgtR0ovHa07JcLGkyGhRFntyfncRrUGVuQHSnvv
LksEGUq6HWKmSrYWg6NeWpRkiITI8vEwK5VKct/jLomHdX/idvi+xQNuE8T4/tLt+5mG7lhpzYyR
p3ChdPoy9rDdNsu7LywwscE3B8OfqebgGRIpU4nz16p5c37xnqanZs9yngHrpMS/GKUYjmWPTEer
Qz/wTAASuCWmC+8jfVgRUxhoL0ftez6vKZcFfcM6Ii214yb+mptoSN3R80AQ0uAUuDndkMRd/7pD
MHvLvpI5RAal9QevqSZr6NBollQJ+QzJGfe4toF4oD+XDiONigZCLrR5a1RlY31YsO0gMdEfxwa0
iJLjBk1MowMs7mqIvioD7UUdg9zgb1I+KiDKC3CgU01zzGFYglxEp20B0C5+djt4E+rMLJFUnOd4
a4Jc8QtLpP8RS8QD8TpX8vKXf0NwKFwg5t7V34Up8sTFQMx/DZiGw15Y8qOKMc9ShRwfIUxH9A0R
iS3HLFnTUmU+0t0COE/XnuUt6l9BVmrCxxysyXfvMywfpRWi5N1Hxl6SagDDtfNDb/nj/nYp3IKZ
jSQKaJukjYcUG4RGO24YYzI/x2xyE3io2StaUFuJIOqI7iMKtrf6dQkqT9nSXZNZtZ/89GQ2pGly
N2Z2ot2Ys2p7E29XvQ7lNbe4ZiQBb8ipvIWXHKGLVQwy9rAHP6nk+5nvad+ZCfc4AzoHZ6VBrG65
b0bKzak/2AUIN7BNn02QrZ6a1SMb0jdZ3Imk13AuJY6DG3o3qxoTJdbsCCh5mu6m6KyBzc3aZ+i/
3PvLy40AKbz6BY2IQcGNKlv+YVChCvSB9hhP001KQoCrzEpEgyf82nEYxpNiSkpiPXMLKVsUwrBq
t1HXEG4xg4fcCRkYLTsjEPasfY9gNwY1mgWL90uTgmq+quJ7HJHS5lVRHebgxsju2MC941smw9Tu
k4VlJlBPs1+9LvhoonCCEYYCSzwCso+ZMxjYjFNjXFXGlbYsDDyNtVbSJY/UoBZnqTHpJZdqu5wj
NS33zcsXp/j3CPEk5eGIh4WC06iASue1xx8rLUpG8LsMzPbtUQ408Gt5yOXS757PVh5hYLVoIriq
4aSIe5WWQDYhfIckHFSflr392r98JBaWNO1Qgd1o0PLqBtWqn1ibEEMA8At0FzWvaN0PUs6MekBH
b37R4eo8yg8N46ELBQuUM5NLlWC4TKHjEGZB+B1vYAwIoJxctmoUcSDf/ZZXnDHK3Vo7e3lcne9e
08DFIh2yB1Mqa/YIOaZbIGzWc3Y9HAe0KK9bTV3p1wXYmcFOxtzPKQ1mb6WqBDaiHnAcBtO7uT9r
MBvHGTCFR52KnPCHVCnpngoFRj4QuiwAsgllYlgzYhjPamYhR6AYoj5HdznsTF0v6wh0xQUpFnvg
qRW26SpwL/L20nhaLXH/LwcewN73xZmluFPIqATTUpL/jy66srZutlx1xl+Vvk3bfoyPAkqWXRIT
OUtWQLCuStSeI+Gyvq+v3cMFeQX/Ir3jlykalCi++inQwZjQ15ta2Xs6hK6Gd2Qu/A/5zBZvvaax
3t/fHv99UUTejvZsisjEQic2JW+zw8s2BYAEovEHUJSQjbXvMl2CckwLv/x522HSl73wVsGDToWS
Y338LPwdcwfFiKSi7EiFYL5bttVinJe7hKQAzqtCKRmQQNzxyU+wl8yrZDXc5zPH+Fbh933BJ6bS
BBLmNQJMLj5BgSuvoOk56ZgQ18WouUfPJkgsWcZkdkJ6A+ggXbFyWc8X5ruarSkzUSCYj0XglsmM
BBv1r34/x2QvG0pdD0+oQ41AD/U4YzD30t3aoG655EcW4u1uvqtH6V7jtBxgqqfF55HZd+QHL78M
HbseU53kQe/mGGvXamJY6sjDEbe9QdqmHH7Zh/8OiemmlEZUJcV9pX30afg+sl0EdjfbdRe3qu6+
PgM6aQ7hqkzvVmuLMMiCtp7/utY03nEJo7eQmqhv5QqOQxHkW/bX0UE3LmIue7tiz5pgfsTzhOK6
lnZqTn+3V2mCjZjjkuyrRa2Fm8I/17+CNBLuCh3rPtDe5TT4K/P2ouuGVQKGva/mYzeeJ+fAg0ep
7FNTfIMh59CziLhM0osQiQWw0zdoJ8T688JU4wKCVgrq4352453FWe2ybVd/z3M8YV96yQYuTiQs
A/yDABnN4nVSTct8j1PnApr7Gf797FGOlMpN3S5BDGfr+n04iLqUabXw2e5SXi7y4HqdxUw/Xssn
Rq/tHN3DqeYDUGozg8EPTg/LwinhtyXJl8M0nj40rkf7rXdQf17ushvIAQGS5y0FJzQ4tkQOITe2
afpZmWUugTb4GYaHZvkPYlu8DAQvPv5tjzxSlEFaNgir8z1ohInrCZXfO02SlfqrkZUFwyIM8M49
I/ltKGUWQ9a7Rm1RC9Svz3AnCfuDQMXKMrL+pcO4wofdHGbDosB8aoJcl0AREI8Jwh5YwnMIVMPR
cuojjA5JHf2aa4vInfkRjj6mkNqbH8Y2+NnDeBPySTyJ933q+is/IlPLHqfI5du0AHOSnm2MU8TA
WJC/jQK5cgquMC453lHuM3MBx/8uVV1HkycobgCj1krlqMmv4M6KMF0xD4IUhXnFcgi/8sbxHleV
JqOqYm1bLfKU7RFFlRKvBAZq8GUR6F/0vTRySmTTe1fMKCqxD4kd203wNrI2sWC0SLMZY9tl2+YN
37hsTr5hEyNprjHhl3taCa4PKZfmRKwb7dhrpNEMFuxbWctPQs2bgs6L42P8CgkyQ6WGJmnqgy4q
bmg6YFpcHpYh5JTFqAZKG+deiLncRMk4XiIl+d9GCITylCGgcwxLv0AuTHAhfFSyB1JEcPXr7jkn
6Th78GqDa1LSNWs91EA2A9sZdaCoF7B7Nzpd7kPW0EYPLiTFKSJIm/AsrRkE3arviXE/CaPvxofm
pE9oSoHXXWQkjli+8w5JlHjErOrgeiJfKumqxo0MJaOY8uOsAJedO1QpgOsia/v8GcmF3eTrJ56V
djZPMk/ZU95OpobwaIiXbu0s+Xqu9BFgAE08bafFtSgvAXnw7Iq0/WoeLOn4AHjzxp/NLBSquc9B
6UF7K95Cl34x4rEbOzTL1PyAPzwXPGh2jlvfUZrqDXd7Dag+vqbZxTNjOBVyLZE5vt6Z0GUavYnR
WwBoP542zbaw72jODWwMRTcfGBWfoLcW9TVdbEfEfOFFFJc/8Ffir6I4YVFFj5PkWP4ihub0PG6v
k6G7hQYQYYFvZosZDaGUE3LPlsYDpZvr3RVId3nZjc5qray/hetjQD2JNy9NMy8rOgSHuxQZQvP7
N+tb4G2KY02CRPBti5rLTiX0inbcGtblBiufdwLiuYBYNmmBbl+Ep5k/RAeHQKtsO6YOeai5AoM8
BKP9T2NH8XJGdpLBDPHVht0wYROgGOPpZek1L5rH6kSLTrAVMSEnqLeDpHdeaKPzsADnQXxf9Vib
dONYpU6qpJuKFmjJgtANOPAFICX51zvdLuRTQWL7FTbTi6taltXOSrVyTJcWdlag4injGDT5SiP0
APLWClXxknuAuuiMNW40zhWHUn4OsYOahZVean5jmUsCMFPuLkyDpcFcDbnzzCWDAy6xYESjPoo3
LEcHXyaDd+Dq3W231VQLbzmDunTnLmvoJYMWGL3rb0aLZL+sPGngIMXXmjx3pSkWQPb+Dt0RTMPb
IpApw9TId2fsomYcNw6/oHC5ZKeW0gvSVNNx5NxwEfP1UkYtPYDLJ1aXJN87g82HkE+raCBRJbdW
HwclEBIJSdceA1yCHnbXiIXo9Aa0lsC6hJUwMuKbp0uLPjmnqOMbhOje8EKl04VyStZGhTHjsQdz
3tA9ZlqWa5eCUMn7dwKCwfrXIbkEwhH3UDlgGMapnvB62inpcaGJEBuTqPOX/KxNlv0YIz2R4ntd
uKLA1e2ygPWzCIYYmp3eOwYNzvR7A0D3TYYhW17FeBxqP43OQIrUEC6zKp2t3la4qG7NIUFr8aT7
UGkqk6Mk0xRVynKV3oqmOC0J6jc2zkP5BInAWPifpHcRW7T6KBOyk25opnYu55ygSre7b3syg4jA
gvVld5l7e3gq0iyN7ubqK9ln89TIQ4N0XrAN7rpzA2jNBcku4sKByeyuOxafF7csAk7CeG+x8ubK
5T8RMUy2Cd7NQV5+Wlmdh3ReaKUExBB7FA22AbK84FkE74C8feX4uBAPnezAduQ/pQUEBb+q8AbY
xfy5cNql5XVuJmDQW0UHFcW9XVwDUMY1bHwj6mn9kKA0/ng9W3eadURQqjSKQJ8xjYhJ+JYysODf
+Bf2G3NdFImYex+lEu07NWXmAtUSEozs2QaMg7SEXRGN848ykiO77+g4Wc7mEp/oP3LagyQGcX2j
gblQ5QBogM6W7+v6dGtvtU9VmHEsSi2qBfo+2m7l8vvdl9dTihx2aA+6zMaisoWb0yhyQ0IH40bX
fvSqSbGtqDhUY9fg8r0YCsuLNH3KuI4n6yuQIUtn7b/Q2kE6w/tCht4KFXgqaFVgfTj52CESlU5F
sEtX1D3bS/l256h37jdPZfV1r5n09lI9oWIsgZh53l23aAmawRPMD/LXYzvGTi1nXurrZns6RRbP
vn2pjke+TpdRXXrb97kIS/M5llQ/0RVGStB4E31DNVDQDUfm4MhCWNY2IvUYVbr26DOB4u4Hrae8
iMaVt8Fr4DpJaWtGNRXoSPhFVLbTdRTGTW69kkmo3yw6yax5anCNYE4JsL2Yg1F+6SUk5zy2RCrz
As254hnKliX6H/r8CgbeeuuB1hafXHKrye0/WB+9yRVEyjWw1fN3e6+V4puIRlxDQpQSseqq1TcB
3IO6oaBxDnAIeEKDFkY//XxiQ6RNFyvQ099ZQhn8yAzj92POToDmdbc3ymcCWlQ49wITr/5ZZrds
DdQYlBfQoOxWQCoCvpj/vzFhGFeVD0E6ss2qXe6mU+5zdAWtfuc24+Keq4dgYeRBdGjaoNM59vHn
omeZAqjOvSFQ0rx9DgHXmFVuc23eRFdAkzsWR7z5uGDVhjwbCqIhUlOedfZOfdPfh45/yhUIdt+0
9mXx0DwCLmSjjimqVxgdn6Kyt0XZoSCLb9rr2UeUgaIq23nk+KcYN+TBjUNYlVq3tDSrJdouaMKf
goiudG3Nfp5TryZnruLRqw0iFKfRfFt+5GDcfLY/E8DB7MStdoJtY5dJjcTYKAQDsoR8n2jsge2c
9K7Ps/Q/Bek0hUO+GolU0Qg0vAyv7KkaenSBtwWkXjGMXlQMqOfEOa0f1wq3ZkXimZtbaxSjgcXa
uKoH8d1l2SZ2oWrQ9mtBpzRhEcrIgoMmbjfTuwj19q7Q2jpAeUxgSZdv1IUDuE7xLdSlYkMDX957
fsDqT+KkuLLvqGR01acmGScVRHlVZLJGwCjEXvQB4yAUUUl/0o/R75fRNzYO+Mds2/CDkA1wPdV2
FOROLjtNbaYcB/2iQsJ4mTWasXxfmfwBOJUFmpkNy1wIXcS4uyQKtx+8EudBsOoed+5qUJAyqg1J
1vlCOva3MZKTHSROOTn6nRkDtbOvuxnyrFUn+ZiuZjLwMeV2he06qGaIS2hRWJvX24+DyCRkd7+X
iErWRW6vV3Mw6n7qt+209Je4jE1Apu9jLWRm7Y/MoCf7LnYbtkHM4INeeITLHSxNMDyoZQX7Lgdn
Wo7/t5xgIlh0JWwYOs2jl7ifYJbxBsAbSLVSlptN2jkf7SII1F80xFoKgIwrh0GdfoTXMuwmRxik
DGfb932K9DK8Oz7QnYsfvNgPzF3zMevRrwreVgJ49ZsWNT/y/2GvL0Mpl1EUzPMmUCCc9GmqJPJ/
jnRcSWWMRkP74B9mYHDiE3tTMeBrUQHtMw1TYmsLtc4Ve7pfDFdeSOCrLSH7hfuoaQsYdlyY56wK
RstOgofB8Mf//kmqbZXoSlGzZr+F4jYukXd7xr20J/gRteptNkRhefcabxjHXqcomTj4twprZzop
b9Z7Dzo6hQTdqSuWp2p6ci/c4j526MAyEBq/bfkgEZiIxxiqBVtf60PlbVHm9kz7KnEVohkym2MK
0npzQDXdc/fn09bEsh4YWJ/IbERud4Eh9eCkI+/1IhkQ8+1JWpQspLG/Mlw7xb5bLPWbdIXkyrsw
Ojx6KaROVUs5i/7Vux9rmBBYqN2p4BdXs4tO9rFFeEVw7oH099O6eYoID69QAKiddqRvuCvcaiVU
nvdmcVgJbFBtPEdqxI/cl1v87Et/RDiVaY3cya1tK3Ioucc5xW5M64T+3SGFvwalZQxynNakYIDf
r6sL3rg22Qjmp7TM2Ek6Jq791V1FQv7qoFOAv51MGOpu0kM8C4psvlI4gWnkyUM5Q9l0ECDR6wfs
mhZ6ulXbTQRub/0BOwUiXRcYxW9Hks/pex3m2THaegY2SFeJUTPIHSmM1cPtd4Poy+5mXSwIsv4R
cGCoXOuiD+hj741d16nVSbIGRdsd+lKsUdXXdf26Nd9Grnx+UY8d6iu8vPQwp+QlDMPUYl3Zk3WE
hFBtMy2AZvfVmZMo/UvA9IOmM0PmOImgkccnkRqkDt32tk05tR4RpAttDYmOau5pnQtYBsC0iEGH
GQCYFX/BNiTjz9tgNJS5Y0AcGNswU7oFjsDvmi5s3LDp0Kg8rycwQylNmgoCCWw4IZDBpb58Wkzw
4pPw01rLBj5QFL7s7JzkL9i/xuR0b7dpt26o6I3iGiYNtlzua92xdjqveVL/mgkKdZXNFRsgbEYq
UkO/57GdIb7n/Lk8AOACDsFQ84gxu2ZvOhD8DYu3xIqvbWPLMc0xQLRsiHYDfKL81CgTQO8j3vTE
NGgUfn0cHFCXIe0G2wqBELDgZmGVeXyC7T8pWHqaTPmOfnI22oswW2JcE0KEqMES+2tQURxfcr50
eTQpynvDQvGso55Ov+vvpLlJ7RAm2RC/p/2tjTp7n3g2ExaJ5yIoLKt2DgFpfAiJlPLDkbvPOK/x
MdDkXwFA/xM1zp5cW+funlIyjH2/IdTWt0lO66/C+5cswWZcuMT0aX8vvU2BMklsape+pkYSoGcH
LSunAHAycizGudNqlqrhLbavgFSrJNLU05yesQysXs6+AdEpRfcJ3C/pkGRYSzP5Bp5q5WKD25hr
oCiZl8S5BipHHHPiSzmrSCAjDsgUx6y6zqX3atnb1c2bZbg5GLdk7AGceaMZ54smejIPS5wGkqE4
7/0uIhe5wD41PiFar9H1wa59AmIbT6XhsB0jNQqHQVf0/gM4KoGKlV+6iJo405Nb8ZzlWRzip73u
OWqkxkjzbkLzRqEz7OSzT0uNurO5nbWB884TlpHTaQoI7RPk49eUZaci6ANNUPgKm0irHAXDRPP3
7rl+GTGZMjTID5qHl6NWCo5y18Fv1AYe0f91igUzrrQnPVsvRCn3+IFIEXSJv/cMcW7knjorYwHx
03qgeFP2iZ5ydL4cixHdgHGUmMda0eoD4GqpzkVSNigcExvxmrnH5WpO0OvnEBk1ZUnB8z0nFF6G
dw9WRMRwq+7dn3ruheH4I9W/AqWdKOQ7YXUYBipzCb6vXb53a2lgTFz3Xkw6/ZtzClEAgKbldhGJ
8ZwE8FaNb3vAFBXL56pHyGmhP+qE9pUl7ZIJhrf41WUolqaD/niLoed+669Joo07wRi16PDf4RFP
lWS/YwoHn3hcSUVDyD3dsbrvUyDgbMabDf8wTfT6jOpo/BFAJBgXuaEpPmzUCeX80Fe6m7bVs9wv
BRBqDnY+Cu7iQnjfsnl61W6r/DVefB+/LiU0Gj2mpwUj6xXEwhUTtwK4UbzvqtzKKqlM5beoKkRT
Lxcsp1T3CJW0Jtpy6VmxbJNtJb/tveH32Ss2Qd9E2ezLwY/e/to1vnx7AcR68Q11IOIMHQ8tioAl
rlov4jwFngPmjreBMAgU7h6BNjYtAkkXJVsoICQbWZfh9EBM6Pc1vawyFbyPJNH7MbDYQ7IWKowR
GhVKe8GhWarK0CLJS9+K2j35c7GhClVCbsWyQKbcjMSN5O6jUEUo4N7zWkT+32zS6Dlaug2SZcl0
+C4uO5Bqg0qqiFi/jReeIy4HjhP/tbbj6LwRI70va07BJl0P0JNSqsYTGteLyt0j8Q1cl56Sihjr
PeHIU/wIWPaHOAi/nCxK5rZt9u71AuWpG5KsqJ4ikXeKnEOEJBSQwMb2azNQyrejdBBk/S5cq0TK
6XloU231ueu1KhpjRa8AU5/gKedihtwfQqDRb9lwkeRp9iauaU7LAPvkigarGHe5pPJt5Tlm4ujc
2uon8/IAWiTy3+1qt/HmDGZe4fgEj43JuGiewG5+1u/eOwTcn+apsF8plruiQ0RRjW/F3DhD2kf9
pnm4eJrT5yoGtU74dMwgvqKz3E07i4PpIO6TNCC7CSb/gNQTPOCSLD6lQu8G2J1xRL2U8U4bo2ey
hyjFZSsojUYvuxi3xkrhBXt4irUtGZexz4q/RdMOeXhvzm4d0jDPShgnxunfFpK2kh33bzOnzly/
f3tgIoVp30vxgVLM/SAsHQrCFQj//sbvIEwfp+xrkd84ERk+9qTgZy8WXUIuMqT4UH4KOI9glD0K
OpM7ccmrwYWZo1kqI0OmJuu95mfjHFHs5iA+p5m2y00NxOuq3N43fB/FCGeMcIji+HhViHjU9a8K
AJdtHZuXXy5KhOhI5PGrgFuhFHRBoQvWJaH2uMP/TQMHQGAGBNPJ2U305fbHpnNQB2tMdAl6ZpSz
wSxNo5YhFnmC/c0gvVYl9n/mccFOiLDIaWvWgmj086u2/COM+lI/+qvqETc8pS+BxDaXgjr+5pFX
UFZGWm1MBvwfaJxSOCUb8j/TL1b6yGWlHjgv1szFJw01s0nBWEyx7myKKYgrQ+XqFqp/UpuBEZYF
D5qa3vNzCACxSfETNb8EL2JqQie5PICdGUHp7HOl7+HMuVVz6Zgkymv0JR/VLC+W54F+HOrhz8fm
+hut/svEUjyDLrT7CLtUV8LOby/rBUY5yecXOhfQ+8TEs9RzIsNOIMmIw2U8d32/Dd4jBaBKndth
njCNZ72dZFk89D2RfX9xVw88aNtdegzdSb9MC17hPuFSh4EpmvfyJCOPPe6Q0aVhBz9C+CUHDIB1
WYjUx5bog6M6srHWBbej66/DjrfCyamfahGP0oq9eRd2zbDc/6O+itSsHvcp3/uaBmEIXef1pXiK
SiBySndGW3aGbBXU9b44tVcOf48f4PP5Yqqnt9wWK/FsGdhHNLOBvFazv6MNm7OWDVX/65Xvcbdj
jJU6UHSi+i7GfOvcB4hYljw3Ca3g4GxPyx7gIG957wfRhsVmNNYTV0I1kHqmw784Qc4XmNnYb/nn
5QZsLoHNl8XQ/N7TMsl8muBfeu2YzA/dQnvboZX/CRoUrEamcZM7SGIac+aB23nZC06Y2BzlMxCs
e7rMdC7dUqjCDGFpMmRMGWxhsEi4yb96MxVy6/K/oZIMmg/Qmq2cKuugqkE/fAnLfSFZe8MdhIJI
XPxcnFUPjyB/HYtggX2H+ev+vz7GuywKFU3XM8bGH0f2ixevCvPVy5IXCRxgwYaclfn4jdyBmHJK
MU5UV3MBypNqApImAR5pipcBnPeM0GmhLg5BnJHU9Wveo+yW03N1I8tnGvWvivagrhE0XXEjN/4N
wQTi/SF5XBsBCgN+ZA2dhOzJ+qB0MjwNQ+5Cu6TN6wZdBuX3hAjIrV6UIkTVWObuT+zGrBDucQzL
BF/UM3kyaVYeY2Jpd36h4RVLJUa3Dl64GX/IQHkgCm0wuJDgMBCgB8SPpHtzm5L40N9RvkA/Oqyt
N5OfbxSd94TxEwrRHy6pABr43+mCS+rV+c087UnQjnygppzF8b8ITxlVOrnLNPKnrq66PYJ2fQYz
YKIt+DJlcxwFqy+4yKOvrVW3HtBf/hwl93TPGSze0bQHqCXxz6v0Bn8CiiBsyQ7F6BKFHSGJLxKk
GlOt8YymIiKowesFG/ACGIF18bcMOXuQQQzCXTjf5uUjWTG7X8tWZwQG/BqeW7801elRS3XvZDdU
gv7Tewu9rqsXnCg0JCz7CcKD8167GyXS6RKEiA0g8eBFmXLHJFYCFce4uwob/GQicpuVh7LzJm+j
A01/wU2xZKnCmCgQItcY19KEYCWbM39rgOB+F+xf2TiwnAp0OF0f6HXEY3dlz1AKUeGjtQOHf3nJ
pKyHhRLnChl+iBKUlzYc3go5d1VhQyt61pAOd3G3SNkot4Os1oL6v+uAzQ2q/5GUKU2KWGFJ+GCb
VFqrl0ra5T/7i6GBl3uP5vlTBhiKMK0Nu87ZBT3OqDptk90b8TjDktsZh/VWB1Qbqqc5O5Jwc3cc
Jth73GDSoS42eBzIYuQGrs3Yoc8t4AGhRKagofdrrykgvoej8P/Gngs9r635UOs90T8yRJm50vKq
u/v8Je48YLG1EydJK8f86JvYo8EwZumXIA/Z8G1bGqqOd4VjTeAqlN8dwCCsrs0jHb1f9A6prsr5
cFYAS7oKUnvmWLUTEm3uwxFQwI562rWd5ueFVbfAWhsXEHAODuvdNVs8p4PkVSsIoDaARjDIakfR
85gyFOdqCb4v3VRsq943BP5K3Z+8zlpZOqVkoq4sxH2yrUgKKZ5nNSCju+IHmwH8x/vZv9cVxVqV
VooT5cEm5QYjoq2Aef0UbxW7EvXbZTXy7+TjwziJhAB5l26dh3B24cL7KvL4njeUJSaUmbFfJtGc
Q+V2zbFOYHMJNaxHfd2kik3mLEgQm3wyuhKeB+Ny4uPAEtfRjQugE9+cjqZPl2ViXrIHKn86ttgP
ux4lyhNgeq1jKY9kFl3EmDZnNocDEGHULgZWmPBmgfvNq6FuLiYYBcqjslnldtbwtdGcRzrFxjnE
JsZltJAiz0VzJlZJJXkHp+qMXGmkKLo79fCnJPCMi6qnTzoJagDduljekIVG/riZXZ2BooQY0cCJ
AtF88fYdDffkwvTU9dkjbEDaSySbZQOAMfepa4f5t1rNdUt6/GTSM5xZEOJ5uiI11f6N9SSx54XX
qjecfodO8Cll8u4GqzC9dvoa3Jc1OeSDpahEB+hChEZB1Nb6NjvW6CuEZwNyBdasLsA4ynOF0cdD
nSVthhiLvmlVcbSDySVFlP4DlgppJcj0sjMJYH5ceSYbicPTK6W1losXdJHQadx/uPxKdPGsU7fL
EeuoaQ8x4XLtPHhtrHOwJdZivI7gHaLwcpY8cpMV6NUYpP9z1LMDIDgiBHXLUQpVXbS+9odYnsp7
X62L28Eg0INwU6f/FoTwBUDz18KjokIUjUUU0neMdL3qO7OY8PRECygvROf2WOE0vfaIUxuPyEiJ
ttwCJhsV5hmxGu5E3skh28Qw2nT2p3nAtYv2GTSv9DY7LDWTFfXHteoH+NfSAuq5nNwo/S1A8x7T
xg13ZalC5pvqUoOcgBWyRxI09vi4vdxn9fuXa6PBjx0zh7ZW8JpY8yT0G38hPFlrWLy3Ed0cH9iW
bp6usYppEJuillYK7JGkD3VfM6U3xzxx7pg0rqUcU2pcqaG2gSy6tlM6YkGq8u8EE4nEKM5ppzh8
0xl1x9ER+fwvPU1NZnIyLDOCIXJrNPIK63VyAced8BRhQ2QRxHfEZLWEXKusTgTbsJyY+pcs0zIk
rOe6qzhvTOrOGuB02flygrNWCwqZp44J6If4ETF/7x6siVLSCSDIgCC9OZ0L1QJakmy7HQIT+P9l
Ytnmy1ADx1sM8LV2g6sSLJ6e9PyZ0YLaoniXOfP1UT9kDHZdYu/ju3A3DbsL8iwCXOTAsnJwFkS/
doKTSR5B4MORru2MpkeYNujvLFqL/Kw4QXkFJCHFq5HYTyqvZ1N99bC2UAevHMYznBeWQbVyLj1u
O/jUg+MblgITyA4ahGXN3XliFO+8fjphuwVDN7VyMss4kkozIAQt80rAYRbQU/uiSH1xHIwYboe/
mZbfRpC/lUPAdDLaLrInVEipnXt8yVzSd85QbdkYiR38BIQlArIJfXE5aVUFDTkpmNrQ37jfcRiG
JW9oHbSxHyaAegek1Udei8Xwk0/miP8YLHUGhbHWYECp6vKZgl+P/QtdnGzBCZFcP/JqOW/oGQ10
pMsuRMcyovLtVXDWSgm1dER1YxGhBbJ/LEwqOMEOQvIc5lZd+PbdOTCdkupBOVCJOXiW0vz+fb2L
VnHNMkR3S+YCaz3pZFtRIvtf/RuquznPplELVap/f5/LzDk0EhW1IaLSdInuajlHSvN/MRlX298O
Xp8nZRT66Cc39/RV3TtVOhLJ1ixM4Mo8WYluxpkKZNORSSpCNqej44ETrYRHpjha0Ijb4tG7tiW/
GmcijpVVNlfe9JYtFSptClI0BBOPwIvGNd0pVvkgW1fNo34WRS4UDnNgVvAX2XsYDllMNZ8AWJ1x
7A4dww1gykSkfcSy5OK1O0LxObVsKYJR7G5G6ah4j4dAOe/5YaP+r7P9RFVGyOra6bopTQ5hD1uN
MBK4m75wuWcRHUAXdYIfUW+OClKChOq1rv6KQiKSz5uzKRdTMNW6VJ38Nb7QBdtECHe97eGAw7yK
IfwRhUctMhHIbgzanbBRXhDQWn3SwE+rLVDJpM2py6eSjU/6Y6ifTFSljULN9o2EOVq9/2oyX+p/
o6rRHy7KA57U5xH/UDe4d11Wr7uozp3AchKouYmSGANwxUmIX91XxoBRxRRyyBrq2know3wXEtmi
TeXTaIq6IkzOGxc+bMusml1UwU5P80fPsRfGG3x6oZq+l217fPZCgftNFpW6+6o6/YKZRgV2U3sO
ijXH4WGYXZWHpiw7isIcS8trvpAyTb4vwoofoNTREVyyJ0i9abvhlD0MVsIFR+UThdnqw5Xh77m3
WQjR/445c4ot3dn/JLEJ+jbd7Zv5oKrb/znhrfG7k3FXsQe9DlTcXX11A2DGma+M/STd2ne60Dtg
lycJ5VGOxrSOHiLbjzRQBf2JukiJaGi2oaS1dJFF8fs81nyyY7wk++eNfxsDyzyzV0YFKT4tOS7v
hYSsmdbq/1DopXR9hx7T19CDH2d5uVTv/6hpvLd5B1vRxYcm8Pgz5UK3X7jF7XqfaNroimctqUtL
69BzDe0PJ9kEAXTy1euMrGsWbJugAQVGJ7CtrgzgKSs3Y6xjFqtVJ6qRmXLRyTu2bWGtwgOJEZ4e
sZB0rwXV18j58pj4DaW/ObjsnB0fHa9AgFB2P/OZyztX6jojf0F500iKLyYIwMBC8c3DQAXH4dDt
0rFPqDWLxP+GnxRtKGz6+46QKEgbJ9BVUhpbSU89g/PZhrzb/tk7t8mV0SvFFGRnZh46l23JMjMO
SLSonHQqFTPx555iHcnvsHrqma2axFVsn6Qfs/hb6J6K598S3gNilH3fLuTH03d6hwEZVRro5zbY
mqtypAEyKDMcJSfYCWdFCWGDXOljfeXG4hdPTCo4Jnff1n0V/UG0xRi9OhjnxxTu/VsuWa4FADO9
3HzI6iZ/ZoxdLCB9bZgo0d+E7FVTJUEsfz5xqnjTtSxemnje2Ha6rEcMNu26SMPEEKcojU2xF1sv
xjNHp93IAmqFDepuQrUP6aAJ3NqWK32vhOfCD/hrIVJAcqZPwZFnJs971cFy0bhb8X9QHxnL5rG9
v6WazJoCcHDDfmjjSoDWEjnKuJoYv3dtVAObVTY+y4V2KNdD6b45r1LW+GF3183ed1CPvSrpJzh4
2Sv5zxpBEdDuBkZTbpJAsGPr+sWAWC5A2k1g+mgbvlrD0+Rp83HlQZ4wtcf0W6Ifmr//9T14uGCh
TA3HZd5v3W3l2aaZdyMrryWtkk8RyjuAaGi/I20livjxSLvlLiE7igv9/z1iK2U+RFACp9zm9+L0
WB9GbkQeMoxXDuaxVzjQcSLY1XAKdP+2maVRnYW5sJxOZRAWARlmSp/cmmFqaDKjq3Hoh2zwt53J
3D0Cs9INJzg+kO7q2t72u5nYT+5RTMgrAviIuZ4G10B36QuaLcbQ9H2h0RDmn2a2LV8xjcei0vAL
8cYjtmnoqg6bGIDBFkpPuQ3yFBagFEWgDFO75at0w5pmhSX4IDW2hJyaVUhSassYa1Wt0BK+9ktA
cN3C8Jx9sCvnzZU4WVCAylN3ux3bi6xclDnb/bRMz4K+q0AB5vEKhRb4IPC7+dmGNf5AScKejBhF
hOaYlH/A8QXbgdVKpEPu0aGW+rropvwlhFvwKJ5Ts7H3h40xTMdPNBnkOkkULcTcnsKWo+xHIiZW
4pYS5acZeQAkWK2Ar7MF8OgFrZ3KF+BiIziEGxZ5CrL+ZsH1HsHzcjGjUdL4jFwjdoywFaWj6QDL
addUFmgna9gOHiXhzFMB8onY0nLkTUin6i7PLpfeVRg2Sam+AyTY/KMEWkhFUqMcQj+4d2xAuTtE
pa8yE0zGDQAqJed41aLBjrpDY4aQdi6r4UGB3RbVhp2Y1qD/xjN6auNiVdH6lElhZFrp/fU2of7b
euYM+ohsbSAmSZg9vUExpvas30gOh7GH5CGmS07GjQcJdDMsoZ8mML8xpvpwS8RPtBQn1AxbYmY7
bn9dvOtpDFHmSvtZ3ATZPFvujcGdFGwZn0drgIiHQn1l1bdI1fPVdYKXtoMo6O/lO4FoQw4zAzvC
mq0jlL5eC9Lk64sNyvEHO0QZSf7kf24B1XjyLpyZEUe/Xm1BiBm65Fwcp6whvavxLgH3YJ42HdZM
sWHNYXKmvHJC9Emc+ZAupL099N98lyjxXVsML5k0KrBeNRfKtCld1H5BME0LqK9ICcMpb9IDZt5q
2H2y2Puqgs8z53HX+X27cmDwbEyI+q0z1EhqSzdh/pejIEjSnRuA4HQssnj0s9mwfaCs5qe6B4rU
5vrOFA6ow5Dq8ByryVHDu2xYs0u1Cx3gAwVw+XzKn4aTodFuXOJKW8kSzG7AI162mXz2+j9cNCc9
Pe1lqNwtnsrKWf9wvvw0ujXrUESFT+Y8Qv9qdQNigyDtQCuUwm2hjTuFeKyNRAE00SSIc3gqg7f7
0j0ItZLzKGGjmat3mSUpS4DxsnxmREUSaHOWU9ESkj6oMg4zYCsbHlYdt3KASz2AbFnl0bFYt/2r
XBKNrrHjRlb/5zqRdnVNcnnwM3bR8t5fGGU3xLDMV3cLqCNcJb+54Z+EEPn5EgYzNdBmfFQrzcDU
Ti2CVuaPIYFcSDMRC0l6AGDpJAlhkCtOC7cQtC/l4LdVd8f1Jztn8qMBYNDmQH9aJw6tdP8mDiR+
8ncx1rJnYvusE86N1g/TJgWXpgli2lql1qOJptlKtQC0Y6KLNyYgtLCrJkGPA5JRsVXkXNvMWxDV
3PDXy+U4Xl72IwqW+ZQ5QKecMVoSsrn/3GOkiyieJ9QsjwqS+GAJbEz0IlHMBSMg3SGwoU/9+zzZ
GhMVrShkh1yh9jzu8mLVN+swKxdsfSJOgxKE3tToUqnWOFd/8Y0reOVpxVUkEWHTJBsT87IEl2ZI
CqXx2PJ2WWp4W0fCUCFfs8jtmcIYe1mGIyx0XCyVec8o5L9x/GvRlTsArpNGa6EhgPiWEA5lzR+F
ri8VrVbZMeFLjR9uBKgUcpZ15Et0Xbl3AaHCICYtmjmkHkYZ3K/ULh3aqGlEeleWnIEN8RPviYXz
EAXCPGWHx2oEPeGmg4nxO1C+/2y3YNeH3Kfs+CYio7RVipy96FMhrBlolA5cPROqOM9Yu/v+sVgX
blZhSx9/iTRPs65dLzbtHzIVIpQuZNoqQVKTLoDsWBc1YBUk524E7PApt6r+5C1WenXTUP0x/R53
zY4umhjJvHtT0xfAO2ROnq9v0gpAgUG0DImUnTEln9yhMWThqkyJ5r63EV8cnVgsu9+yiCygAOvT
nQT+cKFRn2DQOhnrXFHLEblcffqLrcPxMyHFsdgz0Onv0V21wOO/SGcB49LrPCr9axLXd/FyKmyD
4bmluEl+9wtEYi4N/r9LSiW5F97hFyUwGwKjtaDO02heY9Lot+/Ql5PEk7UhQjo0e2sDT45akFew
AUjqad6ojvmF+5/BQP3PSIgYGGH1Vkg85kpZk8MZkQ6LYzYPcYPbqa0mIzN7CaVX+i01SGI7jNQO
hHSSdtvxUpV+8Bkq8+ONY/CHj7aePPEuR7uVTBmw3Ms/Ot5GYMix2F5Z5aKcus4t5Dxhjhk5CmYf
ZEpIgiVSIl+OyIuU2jtpSby/TPk94E4/fl8XkuAD6pwPbRfHBDlreux1SCG37kn+Wc2KPphysY+e
/HGQljBV1x5OHg9lhyqqTWdRBt2P6aOFkoO5V0IXyYypHxIefxLbrckZFTM9lQ/ZY1lBE1SdlU4f
bS4sc49/LvQQcZ2VsgrJzNAZfX9jf+tHbYOmChkW4IyBkV+CLCodjgUrgmSUVFzB+wp1gtElyB5U
cVCj1EliKyEammJign2lUOScXSgoENUEQH8cs29PB3+I0+ExSU6p+KLX0Kaj6YpSS3WOZjBx90Fa
ZJstm40uqMtmSO3RM9vA7TPmDTr/W6kQPX9uUd18ggyA4Pa/tVP16b4QmkZaOredPitYi9xU4WF6
A9Qj1M0wUf+rx0xeJCm6xUMHOtXPSpI2Zk1cHT3Hji6uH/M6A+dZR8vkpjbfUrTFVTY32sbeUOgm
VgISDjlWxilFUdazjoAo8LAfisP0HnQan9WmmBUTPjZ54SdmBYpsSJqiCas25Lez2PMchZ/jltyq
7spIZQFooOzJlMAQ0l+C477CdtQqfWCqdxp+LIakr/3JEt6nVC9ur6Wxs4RAbT4iUmKZ4Sswz5Zi
JURcT3g8c3/gOX0N0ri8ORL7otgGnRJnerAO/o0QVYL3jAqtGSYPAf7UfnhZLMHgn/05Fa4SdezM
0ckW2PI2GLfDtV10gY9xV6o+vsGhFG+WNaSrBi0rZJMJmDGCUnUQ0aK1PMjM8Rr6Q1gAxUQ3bcOA
BoGWfi/jyoq0bE3LytbwXZebvjnlinLTt72LoqSB//sWjtf8Iog/x29cQq3h/Q83EvKiAqUouJGo
mwhAT0hDi9OtL+5p9a3d0AAmEO6BL9IfQ5ter8TL9uQdP83OATIRyE5/h4HIrZfKWF+SlylO5zLj
vsC4KRD0WmSWPH/BPY0+L7AJTjyqWzs49rKVHeqcaBN82gQLdjiSOzMKm6GoXaU/MaAZinDOgmZi
OjdB/tfRT4JGayhIBQHTtfXLT7S6d/fZL670i9cN+1URB0m20yE7yy9feS9M6olDV78cK4sEMqPc
aUrbQXSyG7ecG0tVys/67McOpJkfLcuSmmjFUecn5Hez8JjKpZjIiaUEFgZvEnAdlFoOeRpO6+zv
ScMwZwz8nr0Odv7DaCtyVjDeVntuCBPWEpAOPfLuqy3keSqkLleiVImV6DJTECawpEaebHXV2DgP
7h4mflJGsp6SQar8CanqmQnRSZpVVL39iyr5rT5lGSwCEsdxdGrhbJ2oZ+YvbAhyhkhJIWeII5mp
3TdC/G6BiunTfvDXfI1EmlwKkDvJDAh8RTAIOEHfAQVX2bGw8LfmbEId35DabJpzrLIkoXEktObL
tDtxwGQFrnmpm+mqBDDPApui0xEKyipbgFIwQ3BCu88XkHCM/2dpJFfd6xVC7aBkm6jIDXhEGQk+
/I72PBtFFLQ8Lg0zeeQrji0coq3ID9X3CP31GCemdxIdQUBMfpnvuFxEqowWheeQZR6zXngztPTz
47w5LhBDKT7HRYemd2ljmOgKQhQZfEPv7MVfHxQZ8fCQiGfbG+vdZ7nnY2B1FBU+xSrq8mbPrXll
ovZrHuSfl4jpwrrDBam43J7lnT7VqUv2jrDQ/fBnAsK+twyfKEb7x9dFntrHVXVqD2c/+UUkHWkx
9GIsO85bpGRP/lLkEIBpS5zw+j+e1KlFm9aNy8JnE04rxDclT2OvxxyOVlYz0p3+HOLxkGZdrq04
Ea/JvXDmsg1ciqqCGKPcULDE5DRp+qVV7MAcZ4XtdWVFwLkjml7IKLZroif40CnJT+f/HGvQL1p7
BrHJyEtY9lx1e5Zz8O+5e9ieG7xGmGxdx9Ck9Nq+kokE/j+6PWIGbTYmfy/ToUq9JknBSDmBcQxk
pDtQC03xnsySq1KLMDwJjG9bJfputeWi21cdOO4Y1O3h9z1OKXwcQJpscZnx5WBQE/cCXmmeas5X
bPN7xDRrP6CwrFzQOXW+okdla8/fCrmNFpQUjv8N4pmIGVXMbR7C4TvfQUe9K5r6DoeeFgHkOgBX
agHYWqnU2swlH0Gi84gzd/wI3UcofF+ohblo4k698GGJnQG9OQQq+vYzE6XnJwGBYO4M6kcIIePp
g/AL266xR/xXX1JtlzqgHHB6v//kHQLqydGn2CxPinyl2ZQ7cMOkfr2e9tY27sn3xqcGO62j7NzL
+Ah2nvoHuqVnw8kTpZQBoCK2rzQujiPj2JsKagxPqrhJmZ4kZeycvGl/j13OznPBgSN4+kd+QnGF
VBZZ7Fr7Iihn44PIUCkKrN3SDhHS3E7R0bcSqRpP3yPNpMnHZdMW31BCeJqaZTPyOp2lFrunYcBJ
xBYWN7JKVCbEhoIfFwKpveLQu88HhKPwn6UR1BdKRx5aMBStxJn0mGzsk7Ccr3VVaXWZeeluQW2A
2DWAg560Lz3CVFbnNOzpmwvlLeCwY9Fi/ARlq6iEO4qX0rL+bXzRrHgE35nqyXjvNBRNIOiUIaxA
0j21vx2Qb4kV8ICld/Tuya9jezOd20Y47eRGLCYwtCeQQHkDaU6NWKsb2zamkJ0n7WTqMYJubSit
0M4KYn0g+2PXj1xCtjyM4tfFoha560Ko3jByVGd5FdNjjR0YHjoHQ8Fq5rnb+7h+/C4tWdu7Sn1G
6GPeYLJpiJjBsL7As3Bb7F3r4mWDfwML0XD0TBy5uU9g1tA7hPOCkhCqSvwdULOdtm0CWGOArC+u
JxmSd+2MlsorxXkv7hOBuOOioex2W0zdm9q4D5OBAS0yVqv62+IKxkS2E2wRK81WA6stzECifT/U
s0JCvnc2+oW2K2urDoVXphDrYmc1KzE5w3RzMSBbiyMh5S+aRjNxAGMPbi+YlPT2DIBES0db3cBt
lMhy0A3aasAthVQlrQulCJWqTFkmJUC9OZfHsmDtF2r8T3zlukDPEe/mZdXY10zuOdmHLd2G663p
hwGfh4FJNB6UL7pVdkxxvl1B87+Br6Bra2LGIaXUVF0PEXW+nMn1tBKKJ3h2fIKuCUAasLWs6lV4
oNqGTDS1zN09CTs2wjd4POaS1SXGVi+WkFl6jGqbtjdVgzx49TfNkkfdpgrxa2x5aDFk3Whacnl4
ei11m0nkuQJodaaQr85IyqMGjaY91WLjwPzS5eZ0+La9BpI70Fd9Qd9zg9BA60Am0D4wt4zNdyHO
RPF7qj6Rl02hlCRhfOD3+rajJNsjbseVl3xPtsMm1JXymrwtMVK78uq/HJmUAo/OXOB6B/Jotfw7
A5KHO2unkdelSwzIJVL6PYWUt2+9/tv3sI1TPMnUtyU4K1fwzQXiaPv0CicoUmcIGrQC7oUt3Wzy
rSdw+R5iNDXN1EIY0S8t8EZ+SmsgEIvXFrfW4bwx9PMUu3dkyNgRoFqH0j53DPoZ+cF9h5SGIiNE
MBW3/Y0jG5emMYBXzS0AjkBlXmG2wItCaHm4zgB9EJQ1D10h0wmU0V+Zh3Ueur5hDN5c9aHbCIEX
cxfo8zYGJ0Rj5HpuLlkffIIbiDFVLcq9AwpKqWuAwG5J9iHgKdROpBtDSbHqxw7gFotWHjYXRvRe
qF5zURN6NzgCk/EVYEEG3lW4ZOH2qFQ+Kocz182eGvA1+leFd51aGGQTFc4oHaGrjuvxn3wQcMmu
bJD5ttUO56XJP8Otrs3bDWVFnsm/61sAwdBJEk358m4YxF+TrwF/O1mnvfKJ+7MyMdHNYFOrVKJ9
nsYO39varPIq3MptZD+CcnnfOx79ygjKHCx7/yf5500zhHdbFwt8VzQBGE/VoGmTMV4t9t0HQ4sB
LgOweV2vzLdTjZfAHrAauLcNQZtziqKKT7leDGZyKW5kbxQ8wJgKOr05MS71wgSOCudHDb0mgKUk
M8oynBEeOG3VTa5Z6jWGQbRL1O+2M0UDf9mLITSIldRPSOawVoQwNtpzwe9tnin6U9bFuvQnHrL+
62Lv4GzBjDHyc7RInDFk4/EQIGqc1GtR/yPX1num/16T0kOuDS6fjz3ubUr/0SM0gw8HgsHrF7Zo
aubrrRR2DJq+qE21EndxLNvlvOWYFwxWzwo/dPVpRccgUfRY2xQZBhgD7hbbL9yk2WkpqSHC9uUn
Xxx2pWOSWpd8nVJDkINl8fgtb/VpqcTZO9qMIHjgTL8e40rkKkq5199rJFTrdTraIRkhzlvNDKUr
IlKJW8mfaKd4fBUNcCPS0fDyW9EvCMoUMeGCus9gQ/9H/ZGHB9sAi5+BeKss9Wl6uG+KgwenpWMK
7PUR6fBsjjozgVqDL20PtG841zY2tnoYoCzn0SUkB8l2vwjX/iYdqWm4bSXUzuzGpkNPsdHk2/q7
Z4TMJ3FTb4gw46t0wQqEWyZWxfVxV/9oASirlHrxeRjIGHDQaP2mTe0hStLwJ5gOmM+WHM7SONzi
DcTISgZyas74EEB/e3Pcx6oXF3x4Ab9K3sJS4UfARbgp4ZdFuFJbOZFrKaB1L6ZmNdQZpUVlRfOQ
7z/ewWUSQXQMTM76VqXr5SRRHddtxo30gAR5z9tFeGY3Vfa9F7Y+dYtqkpuKaBY3fMbBnsyJUzXx
jeH9FGgW9v0lpxlTe9Su4T9x1Gm/qYZ4i7RRJ3pPyCqFDkTwWLKVlEwqFYWG5OMC7Wn3P/iHkEoG
IHtoP9GQLHL4uPNWkbD0Io8JxTkGJ7VxiLBMBzyXi495jYJOgCFeXRCj2Rqkd/LzbAk8W29q9HvO
7CV1tWtIqKJznFdWd6rzzTBEthPKPzeUEDlcJVXz622KwPPnxnEvl4/jrsCEULBGT/DOC8i+OENW
BX0mP+csu3vTu0fWcINaS7TBdDPcByyXuUjoBFY0kNUB4M5Tm66cEqhAC2pRDJHyrLBVRsupket/
RG4GIaAcf25StuXATOrPxYnFmuXq+ZKGHg1o2CoNqB5FHNppCpPNHUKHowWW8dywHEcbi5n49D6Z
rO3cyL/yAEvJWMnpy3w7f1C2pfqhgo+khmm+FhIfhomSTP/RY6VjQm8M6KXjYrlyxCsTCqMUWm35
c60Ie0eIBq1WRBIVVCCFROuCvKKUlLfqNnmBOkEtZ75giIWXciB1I0XHhLJnWVUedxB3wuVvxRjD
Kjsb/ziVDHddLsEPYxdaAbkmIF5ndPMkOnh/h82PE7OQvVt540gZd0F+NqEinD2DO0m3bsLSRbcC
J3/uYCp2KM9eEIM1boS/3p0iYRHzpuaRAHzNh4rMJQQ5g8WqAyMQjXwpwSU/hlhn2Vn+OQ29wDww
uVmHavRmETq8l8xBvRRHtBL48+7Wl+/DDCp4hxsgD+P6JshVJMoobDws8tbf3NqwxBPwY4KBx+4S
VrgKhtyjONjGEw+bVNSQ5GEvV3ORolLOREynUtnsU6CYuX4OChU5hcgT6NgC1p10bXtb4/6kUjO7
GRbUindAuf5fjol2iUYpe46/iGPfUZVwgoRjeYTZcEBBn2awuRWNshNqJ5AOTQFEQ6q6E8T/H3yk
G3bCgQHdHHLMJ++Z254XQTXBqMMJkV82Mqck9ZLhhHMn+cIyPgh+05g2G1VfBIn5fGg+K2XcYBRj
whzJz73GJSfhMksUwZVc4Dcl2+At6lPpsxUXtkahbD/MqYPipxrxz7qbpswBxLYjP5GoJXR0ncVo
Fj1EF3VCFQDKajZd9t1KvTwVVf6cUwNj+EaJb6HeFJf0StVBLUx0VHWwHVe8rNOhCjtBvdDuWzrD
aoJa28Cr5tZVlL2GbXZyUkS/00b17SQRLeJPasIe8/6bjJK0VVJBDtYqCY/gzE2u1mlGBBQD7MVH
SXfkr4O9FdupQ0jAIYUhKM8xD56zu3axzzEXDcL9BcAynOcC5dxTJbvU07DQekI2bKGZyPAvyu4e
6JKoe1T99uQ2iyheLJq4rUwmVBwccyJ4IFdfdr0qNshnSOaEFm/lPWLoZ8lqlgaQwBGvUvqSKEIu
G0yx5VtRmKDKmHbS8zxdXuQCYLzfVBKSp3f/2D/e+DXLplM4yVJJlHxcIbKeoGwRHV8Yq4QJ/kYs
i+AoeMfAXGdD3APdu5VJPUhp6AGRiX/NsEjDpzvP+qkDmLtrXrmYAnsFEDPh/Z1OLi7YSvlH4rXJ
HNlHX5tASXOlZ/BX/lGqgMFi/G0EoNL+RI1AGh/3d5h420+Li0375paZsUIxUMFEBS9CYDzV4/nu
vxQEMdc9ksiqjefowcJEnuoISdTZg+zkkVk6LDIaYNJ3gpHqSmWGqx9WxOkyekWEk94fWdM/pzIa
2B/52EncXpz0mw/K2rAri/3YdwrJUUym9kfkSwmIJOX6qdYjpMH7tikhaszvA9zrDWOLcv97D13Y
fxVuWW4k6cgNBfncsKwZ/n/sT8zlKsr5kWQfZW6E2a0rYqf4lkZqhszT57JIfLtXMk1Hw0XBBUB2
K6675VGf7+NMP/j7cJJoO19wyiT4EekfV+N5etlCD8nl2Grv/dQ77GcHuBF6XiTZxkjmehAtKJ7L
gY95C2Bay0wvLNuPYJi758em4XuQOeZCbSpU6R7rMcC0/+7rK28n8iNLh91ptKkWk8/HXGncfMvq
lmNpggKltBggjl21KEY7tecVSuW55B71jP8c5s3NseEaTVsyOaHwR6aCNgr9Qnpl5fv+w9tDiNbR
m/Dz31/UJtZBJjTr1VaYfyBryh9z8VBX8tyamzeqQpJX5YQ9dm61x8qdj/Q4Lnys3MQNSpxtVZMJ
+WEfl4yE31eFWsaS7BMDyaFt66ztQCoPwB/ADp7B/CIGyekiaXmgxTUSlKPlExiqkfpwq9mn9NSv
mHyMGttEtTWqFfYVp1z7SjUZ+uVA3iIemAT05iWHEQD3WW7Uy9QHAMyGOTblrxoCpB9M596jIlDM
t6STPm7gTH0D5pLLTd/T+d5I8hIUwlcvtlioz9cZ3zktFjkLppwatgFfvVnZRhoD7HKzT3n7cYmD
jPEarbmiWtiz3E0ibb8RUG/2S+H+8lzPdfTQIQu7CMe81ajwl8re2Un1zBRmKbbHJLgY7QzRjuSV
hu6OoTf+i15Y/JGY7kkWvKMGqf8U7uNkRwEAmb0rnHru1dnwu787LZaHQSjullYj2Y7QeFVIgZvc
K12/XKE1DbKqJ6RpS9AgEj/QpR+qaGph3VywYCZyvEmbhfxaiVl/qi6o8onf+cnGAQgOtRMNfkAS
2mzgS+VYeCMlbE5Zn1qfvF4cjlkevV/CbVMIFtF+81R7/vBqmA5LQbCDe64dIjDzkii/yjWqztJn
gDzKF4cTiiyPgGVhmUY+8kR/eAYc95CB6B4923Yu+DB4GjkRH93nW7xcjx8IdibctD0RyPaIFjAc
BxWWKb+g3W0FW9npV6dr06zhTSCrM0mgB+tr4FvoYKIVqHZxiR8XfNuecx28UlmFaaE20XZ7OGhb
tITSN4vz71mHtj5BNZ4nfqEayAYYtISBjafaaNrYonNYVFGEIjK8TRKXNueT+iqrJhdTcFXpmjcC
bNji70+ux/nHFEoLRam4jsoveik/1PrIDPhGpCNFxdLMwpzkOC6MIFPZNW8rQ/SJbHZwSOFOw07e
fGB0YaTne/3CC7oc5rz8KeKyWgNDDJBDKZDho8xH8Hi4x8/ylyFgCalXprYKpMa54zJX7SoIesiw
2StTER1LlCtvS0k00htnrn/5C1h6IJ1wPEZNT7O35aOTqPDRuKr5g/EwicQpyPtpaEjmpWLtQikr
hGwqLPtg+bSeOezqmkkfAYN1x1DpPilUJzrJ4TYe9vdpJnsoVIUyr3pJ6m2aQ53WT1vrxglt6LNE
THdbAE7ii/47Nq+7VeMn1bydXWj2qhYDZSCSVcZD/0hKlY1Sru4+Vg1wPrZETt3MpkXo/biyoKiV
hJctV8vrXUnmoEI1VL0Etg+QvecSahWQ7AJ/Ey7giUgiW4KNbgWsWEr2f50gAcZrHAgIWtawaw5D
kSsUiszoocZTngK/7guAzvsd5dK6f7uv8W1Wne9JxWDth/aE3XMnNdEXozhl1kmF2cVmroeBs5mh
qPz0FhbMkP3lM589EYuPFaqnKRSG5nhl0d7SBHzqvJOYmBpy332sFtn8cSzi+iF1S17czGoKKK+s
qo1jBbdnHyGIxXQgzBjVpNbYIJ7p8xZBg0fUN+oYV6TlAqQGy7DjspvOUjiPl51yfKoTVdy5GL/q
hsyTnwnZpGuNk8jh5Zln81ytvD9/az7siTERrDys+y67c7eQ3sm8GovKLFuJ7KgDWygzUd7JxRfn
lOucs8lGBFyhSm7CD9EzUhB+vc9Bi+qKh13yMUr6aAIrD3kh5R8FmUpjDz0AB65R/R6jCc2sdqi6
x43zGIv3/d/0NDpwJKYqhiGVSThxbaGIAvFESJKd4e9D6WtoVPRw4KV3DY4TqeeR52mmVeRrIkmJ
bi5MqRM29UmuL8BGt2wBLoK6Rep6jzNdz4BI+CguytQIOjwQBkqeTxpSDx56PN4ob4GefnA2DQRx
EGWBHSCiv6vbLk0HLYJW3eFlbSCr3kybbYdlTRQm96TmnY9Joc2om01JaVKWjcNpMbEGPqQwar9e
9KAb882sn+KAEx4rYrkOOnozOc1UylLBpWYYzWgxe3yx59lyZ5Hjcni1ExWV4Je2dPCn1pIlpONo
0ycvmR8jgLy6Uy63B0s/D43jzCD5rRXG7YSfKWNXIOw1r+VW5iw08BZndsTwhixJvKaHqIwRWtbo
+jPja7TPyUHN0FLIX/pwF/imGXTTFChUAfmkI243j9rFxfQ3Twm4qYhUdYc0nAyoHQfitRXMNeP+
xUF1wrJ5vzEGdM5+0xfawFrFu+5UDFUv3huMQ1yhmhWikDb97JAEnU3802cMWUjz7TjZYs9BWOhy
GE83Jmyzo7Cc8VsF/Zmiffa7I4pi+uBhlsfFE+DFg3j3U8H7ld4bxWIZop8eKlm4sYd7nGm01Qy7
vpl7ABuHzJznr+dwf0RK2Ui5R593MSJxXnlzga/F5rsxDyflAA1fWUGoiCzsiaT9MPy+ZcRn9mbx
oGuk3GAtZchP25x+X08W1rB2wza/DDv8JkWPHWReS3H9VPSka+2vsKc0kPy+hna1c0CzHKcK6CH6
3d2TsZYkKx3DG5AnBULeZIStVFGDNbky9aHgDcq5MKZDTVAU7rGHEMa2C/figzuZ//HcUcq/RDgI
jQEWR4PQKDpCqoH9VZKla5Fw44UWlgj6iaNE6A7ooLD/pQp0dWoPWYp6XStlw0PuCEiR+MWArb1z
vUU4hWT7ZUxoBn8C31rONPWTzJNgzX12trfmZApKHAACrOh9yy/mVoXoLB0PtLORkwJuv8jJorgA
mpujzuodRozuTGfsERoD5jn3MlAw7EAEstCpCPQN1yvD+eW7WWguatGjnpE8M4qeX3MAniPNsmE7
Cw4HGx/zBq9XI05oiJkvPWjjfQ/KWbclFuOXjeqdqqrdshxomi6wlfyantQo8uzfXZeKvuQbYF+P
azMyI23uV8LZcFvK4o8pwhRLLWRFIg4D3WK9ST9pie/KNSyj024bBtNZbSyNPfWmvnZ/YL9L9S/O
8ynOmvXgTPdUbChv8d3CjaSN/LndYpfWzarXSR1xgIxFn6d9EMSiIIbEGx8/fASd06P9idJlAyGG
+bw42pdQ2Mb9agQyl7nUsprZMGcDY7Y6JzDx6uCoeu2SiQihyS9Wnxmh5H0C3kU905t6ulf7TTl8
8PsXMFqiMzrmB8XA4aiS78WAYAW+jinevUMhC2XY/KK4YyAgKYsAsxrGEgXCOHe+ma4azxSmGccx
gH0Ba1ZjwVDQmXkrMS6F4Gs/Zs57k/OHfBeGHgsaR+fRcGyFXXqZZxdrKVAVlKzP/FJhNJmHhgke
MwBoCBMTfdazUXMbealT8zAsVM0LNAKLthZbr+/j4gq6ay/5myK0MSCfaeBBQMULB/45qx07MD2V
zCXkBhowLNBpg/V7LHbRXHWB5cBrAYyUrOcC1ta2/7hbGK9IXtiUobPWL6xBUeN3bB1sUUexF4oz
Us1rP9yny6hlBOKBxPGWEdJNklTqqp/Ocul9R6SM0Uoz/37Lm4D6KDGQQm8pdajLQ9HrNZx7ddID
YQ9wxhyoLGfRE3xlhug08r6enWvTO/5imBrCVtHeDfW05cSfP1wYCrACGYr/wpV/G+hN7QNS/z5K
bHyUNmyrmiCkdlOpgbHlFHHzjVj3Tn1V0wfdaj9wwKDJg2m5pWIaHQk1pxQ9HJo9npsM/TO0N34N
ORFqLNjhAy4Ovs/B0ypnG9ojdMFjtguhg+LY0heTL5T3ncfnOOfionigC5yQLcZTBAJ27WhzPKJe
gV4kvUrQaRLsMc4taUr4uCLUxrtWJMR2UnFAb94boJL0EYEf+hyJbVeW8Nt54+sFv7kgbdruS09w
IUzbb6Iux6WMPPdK4xQpGpc9PrEYdOUxJo1oK1tOgoTtMwA6ygSnTvWOiCvyT88hsX7iVKNsasR0
P2n0LLh3XWiYgD9tqJ48jYB0s7ykFD8vDr78Mzjo4cx9Zc0EcVeymF5zi5g8kZzQMNQEFkkxZc2l
l3rH6v5IJT+4iAlO7Vl55YK584xkg2BM/iMKeuCLFcVjK4Y8XoCh4USfLnprHh64NxuiAvMrk8/u
jFVRmARys/Tx+sNZeq8jDmdH9riqpGc/w+TuGGrPMguGhi4uiKyeWbzrxZVCefwX9h2Rm+OR7atX
JiGTkluqpQuPg5GcHYRTIxUnEeN+ICt3KA1JkqeBX/BzYwfGjp102KeNbatbVbyGav57BDx9q3Hx
6ZlARgtQFzNR2oR2XyVWGweBP9dU67GbF6EIYwxUKovmtvh1hTQ5zWza6u6JRiu5qaOJ1Bp6tl+G
02sfE4sXWH9eoWgCpIaUSpmdz8cDgzoLT2CDp13jXs9M/WeAVsDH4DJcjH0NZlGJo2Zmaj5HK0Z9
qsoJBiIQCQZw

`protect end_protected

