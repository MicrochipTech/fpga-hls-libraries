--=================================================================================================
-- File Name                           : VGA_Controller_SHLS.vhd
-- Description                         : Supporting both Native mode and AXI4 Stream mode
-- Targeted device                     : Microsemi-SoC
-- Author                              : India Solutions Team
--
-- COPYRIGHT 2021 BY MICROSEMI
-- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS FROM MICROSEMI
-- CORP. IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM MICROSEMI FOR USE OF THIS
-- FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND NO BACK-UP OF THE FILE SHOULD BE MADE.
--
--=================================================================================================
--=================================================================================================
-- Libraries
--=================================================================================================
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
--=================================================================================================
-- VGA_Controller_SHLS entity declaration
--=================================================================================================                                                                                                                          
entity VGA_Controller_SHLS is
  generic(
-- Generic List
    -- Video format selection
    g_VIDEO_FORMAT : integer := 1;  -- 0 -> 1280x720 1 -> 1920x1080 2-> 3840x2160 3-> 640x360

    g_PIXELS_PER_CLK : integer := 1;

    G_FORMAT : integer := 0;  --  0= VGA_Controller_SHLS and 1= VGA_Controller_SHLS with AXI       

    --Added for AXIS_Video
    g_FIFO_WIDTHAD :integer := 3 -- FIFO address width
    );
  port (
-- Port List
    -------------------------------------------------------------------------------------------------------------------------------
    --Added for AXIS_Video
    --begin
    --start of frame
    SOF : in std_logic;

    --End of line
    EOL : in std_logic;

    --Pop FIFO (used to pop FIFO during the alignment phase)
    POP_FIFO : out std_logic;

    --number of words in FIFO
    FIFO_FILL_LVL : in std_logic_vector(g_FIFO_WIDTHAD downto 0);

    --FIFO almost empty
    FIFO_AE : in std_logic;

    --AXI Tvalid
    AXI_VALID : in std_logic;

   
    --end
    ------------------------------------------------------------------------------------------------------------------------------
    
    -- System reset
    RESETN_I : in std_logic;

    -- System clock
    SYS_CLK_I : in std_logic;

    -- Specifies enable
    ENABLE_I : in std_logic;

    -- enable external syncing
    ENABLE_EXT_SYNC_I : in std_logic;

    -- external sync reference signal
    -- EXT_SYNC_SIGNAL_I : in std_logic;

    -- Specifies the valid control signal
    TVALID_I : in std_logic;

    TREADY_O : out std_logic;
    -- Active horizontal sync pulse
    H_SYNC_O : out std_logic;

    -- Active vertical sync pulse
    V_SYNC_O : out std_logic;

    -- Data trigger
    DATA_TRIGGER_O : out std_logic;

    -- Frame end
    FRAME_END_O : out std_logic;

    -- Data Enable
    DATA_ENABLE_O : out std_logic;

    V_ACTIVE_O : out std_logic;

    --Horizontal Resolution
    H_RES_O : out std_logic_vector(15 downto 0);

    TDATA_O : out std_logic_vector(7 downto 0);

    TSTRB_O : out std_logic_vector(2 downto 0);

    TKEEP_O : out std_logic_vector(2 downto 0);
    TUSER_O : out std_logic_vector(3 downto 0);

    TLAST_O : out std_logic;

    -- Specifies the valid control signal
    TVALID_O : out std_logic

    );
end VGA_Controller_SHLS;

`protect begin_protected
`protect version=1
`protect author="Alireza Mellat", author_info="Software Engineer - Microchip"
`protect encrypt_agent="encryptP1735.pl", encrypt_agent_info="Synplify encryption scripts"

`protect key_keyowner="Synplicity", key_keyname="SYNP05_001", key_method="rsa"
`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_block
TJQZ+3LPTirZMtCRG7iQWNGNZPy8efWPEfySnzkwi7FeGljUaDc5pMEngNxa6fmbJjKz10NvX90B
eDNWHZTtIczt79wc07oQ4yCNrK3oH214hZwtnqnXM3C/DLlFP6KW/WiK1qDebYl5wqalYRtoN0K6
cs8ZL5ZrNwuZNbP5M0BAH+AZSMFwzm3yC1yX4OVZSRyinFe1PiV4AnSuAwvNOREegK/e+czuCy4v
vp0Hhv6NANM3BgVhlYfQzj0lfvHn5PS4WPFA0/VVHrHGE2VdPZLocHaSP6Bumnjl3QJS3xzboVe+
N5RD+EGUuB2umGe73hHEHNVMe8/+NMYHq006MQ==

`protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`protect encoding=(enctype="base64", line_length=76, bytes=128)
`protect key_block
YC9nSoON9VwlU5UsErA7RNH2ZeN38ye6G0kevVZcqnZabKER6Og4rbG9JEMz9RfhQyBguSsWxy+/
6ePOJTY2Si+UDEC3xQLZcXPhcMItC4miVTu4QIQ87odQm69NmO0sFBq+yczmeixw8k6q9Y+9YhsY
LSwKOUHPZulPEYf72hU=

`protect key_keyowner="Microsemi Corporation", key_keyname="MSC-IP-KEY-RSA", key_method="rsa"
`protect encoding=(enctype="base64", line_length=76, bytes=960)
`protect key_block
tdJRuEg8h+zFo/wfwtWFIhDag3j/mLW5EQU1CFcBGVRX8QLUdeKRR5XkwWCV/Q49cKiQ1LPcOBeg
jDIcYqjHQup5r1/vA1vHsjn400BXoUAP62XUkxsUaBWWSFsy3pCNaFH9v5aeEuC8unpq8OM37S3M
ggFrmCm0BeoJukXMEtRdM411qpHaA8+pk2ciPhPQb9N+Z9hkHAzcod7/toKc2Tk/jTVvCmntstew
q44CDEq22c1iKqUNPYlJe/fcJyIU/KSP2SPfr0T/5f2zUBa6UrvHlhPuiNtdadiMrtRMTrE4bQ1h
qZesBfcCqyk2iQGQdMqIfZ6l8W56PpR2ThysTDhgMWKm1EkYKWbw7zFrVHGQKJxgnihdjSXoPYY0
ty/1qKmRrK4d6G5H5Ag+NZgB928/hgijgi9xOnZ644i7V1GFinwBD0hxAdpTqJ6Io3N52L1mKwUT
7LFFT4CZO2V7WVyJUvjqlqkQVRMlgtw+H7CrcB1JpdAltAfVmRyssG+M4iSiroDwzuMFw5pDIfD9
2ZOCyy4anaV3irMp53pqwMLb5fcWMY6ZsIj+VGEuE2wdX9eaO+aBRUnc4N9ny4jsuxyy562YexKP
7ClbwUAvFiEw9qnaw3QmY5npqo8EPpxIWeJdeYhzWPuDXNBsMYHPajwn9L6nm62utmei3rlPdNMk
leOE6pK+vXKAN1Bk1lcmTFxu5Yxm+5rTJf6HrHzPFYwBOZklBLaJcamR382XddKU4WrFVdtitcNg
VNLOhXYar5iVQg21CgF8rhe0ZGsESxLMue/B4gIHbKANba9QBZ+MrAjzVzcEN8YDdTeNwUrErS8Z
K0A92hOP2q3yETE4slHQh7LFNAY+CmihZDiFnX1EDSyiZxEMX6p8k2fGWaosUBgNhRJqdhSyQcXV
6cHJrQ1lfqF6eqXRYzWEP8XhPtO8jB5wrHiSez71E+MBBdecTNnookI6QOEUyolCeUVyrzpO+UVJ
dqR1X2y9QLjbo1olIdpdSyFf/53A8mPRqlb2WsVviMebmDPXFZxOyzzS1ej7m0/TyDzVy++6lIOG
Vu0CwTQOUieu7VrHQnRHVs9rfkzz9w1H8XeZmsObkge9b6FOCNdu/vptmZfMxqk5I6jH8pceHwjG
5w+yDiPa1doozomWKQCDnl0o8mmbbnhSCnvQUp3+n+AyPhpJZweSH4px9Vx4GHYyT7rKYkPGCliW
DXnGVKAsFOeifRJw3H0wtqmFHV07X9V1vsZrQGE/frW7eqz+phSVix7cfHNNMESI

`protect data_keyowner="ip-vendor-a", data_keyname="fpga-ip", data_method="aes128-cbc"
`protect encoding=(enctype="base64", line_length=76, bytes=38944)
`protect data_block
biHuFEkPV9RCY82LEfk0eCFMtAUGsK4JlRZsqE6wL0x+Gyso531Zw+NZm48TEgYJeQpxaDTKP8rT
LdDR0xuA0juPzVSuQ18SJcCrzuOkozsnepFd36DKwJoUXiiMYVcuYRj4rvskB1kxtGEhfV+ZTviE
Wz6fyBR6772nOuB/VHj19xZWV+aJ1P7GiY4ifSF5BI3CWlNqCUZl6YRgZmgxtcgm17fvZ0BlKafs
5nAZr3Eh+RbbjLmr9yY5ImjVSH3D8CUgAic19zaeRHMNBwCRvx9CMr1g0Ydk5bLunLq8/tUMvzqn
3LPD1mVY+uk+n2OEopid7gFtzocWYYvHYfKXPNAVCCu4O1B+hp1HtGPkBPs6VbSO2SJhYUBVfpEY
v6UDd58kgzIYS+4J88TUcs2U+tw3+F9vzVuCTiXjVz30uzdsI4KjsmYAlyh9xFxquUIdcYZdgmGr
ETN15E6/Nv9Ml0pez0S8wReG1LB4G4L7u3qkmrk3azitlHC5oH+5v0ubRXQSx5NrGY4QcS54ipsO
7SWW74LZp5SFWZGtrNGNyc9dI1WAES1tnHCRIpQJb81SEzgBfS8p3g08FatueXt/iR5u8/lNXgb/
4tXBzZxOws13xYcAjUcLzCBZ9OZZ2sGsvPK+SC13pmflQaHa8O0Ci3wacCKk5jwEMNQEICuZxdSm
GXts3wmaS8vfOV5iAsm+Cy8B8edQie+Inb+mhrSqfEIz1SMOdnIzIUq8sroZiOW7Zn3rCWHJVpp/
y2ZOpb1qUPmsQtyd0EOyT5deKnirJjLX7NWXBsm3V0OFay4AD0Eaj0SbatOHmhyJke1HEpnmbg17
D6KUGmDeayN4CG8xlUwxecw2tr/0DoxcWWaUgTjwT+iP5GhEr7Xm9RUHMaoYWY/3i1Bj1wgSP8H5
LKVnbp4WuO904MhYIwLToMKzcOjkc/q6KwsxD6t24l8zz4krY4VKo0eZweu8KucLHptg8FKCOwrK
1Jb1h64gA36e0roSqLPHBww5xTslCLEZpVKo0JMW5O17bAAtggMTJQaA/QQfdmEyww4poxnfkWBJ
yHZFWjXRXwtIZ/nqX8xaW8Y7i87CdifrED3lXZiJG/MYSjeirHwYFb76iEj5VDot+A1WabKNRhNR
jBoDnzkH9oiZ031aw/xe8yZOMgV/96uRf0dPUVU9/KY97ZY81Th+pb2QvBx0hN0z2+p/IbGy0RH/
6UtUB2e8xKc//j48zOOs2Wm6XSjH1koKMMtHtI9byYjB8vuW+0cKX8e9JnJBIJHRAncYJCDR5X+J
MnFP15fKHJAr837pNLvKqTvtSG33NlA3WD4sSdl38TTLmNVxtdz0WQMkau28nUN0TE1j7ovuTz0N
haKEu/bpP+TgbR/3I+AamBOXGoU+IeMcHXJIgcoiNP/m+kyFBk6UeMsNMaAzemp3Uq7va7nv12Bx
2LTzgNyBeukaJzczAKXtm4AdIc8s55NLVcXiqIHX6N4LkJANitOw7Opoavcv0HkVxvwRK/HzTVKM
2o0Icj6hJBrwvjTNIOcpMk+foMMAj06qiVlmhlwQmhii/XJSn4fIJfD0Oni7N45jeHLRc50Q8Dqn
sr7Vh2YpwzkctUG2Y9rrmpEgN2MLsN4jcib3GcN4coL59sYtxG5fQcqJKXwlcvEfpZBl84RDBsoQ
xFlEzPHtYjyazGcESniv6hLY55+Y3J5InEuZ40Xh52ysKO9KWYASO1OTf8+XKvy9rEHhmpEReoMa
4mOJLDRaFgA+tIb8pC1T8xH6dIZGUbp/PfEKz3dyQXrYJGni1DJsF+cDaAKSV/VBoKPEgB82wTsn
zr2tt35ChaSSJkeEuON3vkcxkdbpRDww5KZq4nv0/ZnQstl2NiF33fgyuKXw1JYgXsCRvWvWymGh
nDicRqTQNLTVG97o/vD+38uFuJAKZjihkGE+VFHkYNK0MeLWN/4TRKfRzqo5NQcUXbnWQiRSJf6Y
D/S+AbtvnOWu+WCK1nT292SUC8tVwuX2+RaEAmZh8oVJ97mCDVJ3Q8N6/F7szawEnpQwUwbbp8RP
j0DZEel1ftw6QPB4uVZ3nqBNmC5R1mfJCx8YByc+1DPvHwex+MgRc8b9zzAmNnOML6SJoeGH5S5h
82AN6CmBwkeJofS6uOlB4G5emgvSl0rJ7yzbqDcl9yXGpofZ1Wsv/nYJcextOvwJFlGnKPZWqu+8
05lA1KJsfiAN2wH+C+w3Agq0tcG38NJmECO6lJtYa/BrnrteaZlRc91Ox4XORP/lx0/V9+I4CGqi
IpHm/cF0sGfh5UJ8eQK58JxuEXxVnYarQ6nbkO5k6cbaXAg21kUgsxEJpCUyiAF0vNswewnxgJJ6
ITm77W1hjFjkLMJHxGdb1USV0inCkVzDU/pP10tRU5rvCUEKMP+LcD+LvM+598Lj3G6ahiqtz7S1
Z5J7xP/+tQbE9+HoYaEqM6OPE0xm+KGNK6+4DAjUy7nayzAwqXCIL3BnsCVXYgqXu3NZwzb5i8B1
AFgYHCWTkT4nICt1Fk5+p2FJGPKy/LoI/aMOC74izMnjEEEEfhToIPFUMyRGNJyHonp+FpxDX8fS
BO8ThKWgyzVf3gfCK2AclCFf2CTuu2dw9V+A4yGY3qnT7UZEvJmEo62h/ocTkulHtpz6klhHigsF
7nAkBq3u0DXQFYPbDPsXltV2ciWjfyp9w8wdYCJFu+VSsjBU9JQkiItg1HCtIXd8vTyyWUxCRrTW
MKUtRHn+0voXSCoEcl3OhzOtXv/qye5JQ2GZJ6ZBbFF2DpwUkil50gby8ZNbtCHhXduY6F1ViI8m
0vdp8UlvcCOKE5NQVqVv9NVgHevVz2Y5RH1AYVFz0hma+J5DZrCWXSqL6mTIdwZagfch77/fD78E
LHRBTB6WPrMMqQ8Pes/l4yxHUVJWFNJoS04rOcRQDt3dGcCZeqeKwZFCFI2uj61+h4WdEZfdpwN2
Bgy46KGEDrFQGmEWyiABOf6xbZf2u+7mbm1C5EzWyTtWUFTxPhov8Qh5qzMQuo7ZVoBwpu6fMXFL
A6A9mXOevg+fhVKkFDYWtMc0nwIlgBNhztYYo1Uttrgjs9RZN9/7D6UpKpPEJSWQC+AhKe8bLkpK
BPbI9cN0VfHd6B77xfXsKy0eSlAvgRGzCRC+1kSNYytxuko+ssxHkkwzD+CUU/yWI+GfYUI5UrG9
1CKumc/mEa9JHIpaewpPhI0pPiVnNino/XjngRCggwOj6pJe/uDYy0zqqS9zg8S5YKTN5v5LZdPh
MFbJQI4qkZ5BSXk7zOXLJsp26SKXtSMnmWe4IMZUhFbgR5zorIqa5r6l6hnQ4hrGAFnHeczK52PB
D540gIKGbuGeFcX3J7EN/ilaSaaT4bg6E1l7uZSZi4t4Wmf/5ggOmK3chux8f9UQF1KSpsyQW5mL
NbU9BWXGmb7eABmvb8jRpE1KZ5vakZaoHEjnY7o0Q7Ig/bDONamMWHjETaBmcfPRtza8GF8HUjQi
F2ezE5aYDsNY+F1inJp2PJ07zoEvZcGgf1I3r+cN035aHOlMH8Fl83531bP6Er01hwkiUHpu20n5
JBpU41QRtUxQ9w27NkbTo0hwx02p+0KqOoedE/FnRJ1cNkNr2KPr3pVsO0nFKLsEjYfXBFsOU1GP
a9Mc2Lg3YJOnvkuEy0Ba2B8z+FjQmK7ai0qF4xAPSpjjlRjxJ/eRq/RHMKlpdI107g2hdJtbzvWL
KTmjtg/Sqf2yaItMeboCTbdSDKWb0DHLPHOcky3EhKV7rebVd5/RPOHxymDLfou843iv/1nvsw0m
j3ibGmLx0oCC2IJCnCjFqqm3lTz11xE5T8KByDmkCatN/BFtmdEo8TAi1CMjlgw9ZcaGimE3a8Jk
YLAQ6EHGA7/sUd7iW06bIHxGKum2bDvZVMsJd5ApbT6W+N9ZXkAxrGB/NW1BnvaDd2k/2dwpCYQw
me6769ke/c2DFYUNiB2snJsy45r/gMFaph+j2JyLxAb5J+JKdRIv9KHM9jK1VdgLzy71nqnDhR/4
wE80pN48deEbNhKqbHHoq1Rh4h2NfQ96knMhMe5rKXQdnDYq6t+6S71s4KQ5kqMvW+fcsqEFY3SD
dxS4Qr1QBo9PRgG9/ZhxMBt9WLHJnMwRWLkyk+nOjKJzBAN46PlszsbhAapAjstFcxdjO5y0RCqb
U0IArl/dcZxDXG6oCRPlEcYKQVMvXrFO5VH8TNUeMH5MOCwGqgOBP+TZ4G/R7NSfenCeaWEK4by9
ltekbtc/UQraCEfrleGJxcY0Ym7jOCW1QEpPL+4HezzWrPI/JlfMNM75ubb7PMqN5rawm4dsTx9D
VlGfE5YKgrpXUM2SO+jwMVmxbUw/ryusygjIJ2et2zjFg8o/aycjQtNKzOO0KWZpbv9hW8j7sWCU
PErGPeWDW+NndGcL6mtHAMRNxpZoryQX5mC7kqafsxHbwBGlZVtwKZq1sQftsrvXoDE+q0qD1DFc
XZLkMIQwhMhupmnJ5CbB7rH+3h9sfyJZmZwrEZVekzp5njh+ZnmFIWOoQdMfkpaj9Ox+GDVsJI6B
tuYemtNvmqHZUQr7IFJyuHETxYOzfroIZC0S7ehL56Vf9IPRxOsiKRHUOh4jqzX0CuUtB8hdOfam
oUg+ZlK5p+1/8gYRJ0XWTbFJ4T6d94mSyhetag27akzTwx2+3utdpoKkZ6DbrLu8olPoSyyywknN
oeSrvCedCtLfu0Rxhw70k64meqeIHUL+MA4LteVWqZu/wG2v9KM/49bdBir1BokRJ/tNyxJ4kpbV
agmovgZIZXXEuyy/VS0fLwuHXojE+utCgteyCmontZIK2uPb6paGBKerme7Dt2LAvuAmo9SAp0N8
3du1GF4roMMHusGsHNAvBfcMV5cl2GvCBzMbZAdJhSSif0HmXeveS2mIHKYpPtBtTgwM9YVtWFZx
1Gr2jji0fYkhB2Qsmd9uJnJ9hvHXT8detMGCQIPNT1ZQgq9Kiis20XDVEKe4juhm5HmTsSoY6tVo
nY1wOf9QW/sxiGsgN+HypVrSQ9kCSiK+f5miHcRu/2lDfsCB5VoVpKlZeHReUWgqtsEFKjIEPcow
61I3m7GOf+lh4MlT7YcDIj38pYbsuC7AY3S+p+rL5G+g6EEdM1nEP9jZCiPInzilK9HTGfkF0Y5s
vdbaqI7lz9EW0H7p8mNbNSHrXSvuNgMy7vX+3WXH2SatsZXUxfB+padub6qyP9IG1v93Se8A4bOU
SscSjCGKvhGSYjDcBH8GHPhcgQghKNEEZUhn9u24iV7okqQ2L7lxWUl+jBeB6Vu6Vq1JCLQ8z1It
5VEPsn528RtRWpvzir4z3xXlKlmv51W8ZELh9jEeiaqeyySfL8KTFAVALQYZ+MHKCt/Jp5IQ74dA
BqvKldRETy24NnK09iF4VeXtqQFnVmNS/i6cjVrPzl4Cm6+9JWZ0ne/NKH7TJX7RPfv0u0pMJntP
i2PkyJ+M1jc6937cD7ot5DJUpVMpwrgakTtST2gVKvGF7BTQpyrVqZlNo+RifLlWdq/VzXkNUqH4
SIwbdhujrSp81VBBYGahkl86Baj1Lyno+NqPfScqMsGtbjFCpbNzZsYCl6haIzAWCyKPQa8hP1Sz
+ryiG/rAuqmAj5jhgH5aOdgZAmTh1+zQTmAyxhXZJGF9A+C6p6LpBrB3yxpJMLZS/UwRpgQkVUMF
lsbwUFVyEg17ae1fNC+F+m6Tih+pGbcxv965nNp8QLDCpOxIgOQkPp/MEhGgDRuz4jal6TYilHk5
Vat7kseqaRPRJR1OEcEHApUkAthOjNmZ29I0axDD/PzGssF8x3ZDfRV8lkBq3PYSasPTbrlCUFls
QNe44GHYUytPdS0OegF6dUGib95sOL1dPApdjcxOQMyY2MkcQ6uTdq8cJEpB2kGmC39JTc1tW10T
Rs2Q6mkXM0IUfieOTTLIo9wVhvXeCsjL6WAZWkG119wuSDITVM14td9gjz67a9ejoSVPWHjGHS+R
xWgu58fowa9I2TzzTEvLmwnN6vIq9u695GsG1FMPzY8JzwP3gblhouXWP6rcOEGBZHzq4jxTKhIv
Pqu45HZlZ42wywEfGwtjfHl/22a3Nvn8Gh5mqXTYz8e/Vex9eZc8x6dv3CDspVNQcc90d0VmnyHK
6GZh3Plao4JxmIscVc18Fy3innC1l7ySaId664vJypbwK9S8IOBoRRfjtesiplL1phNgqzHHXJmX
gwZH9InhGGotRSPQ8d8RptkcJv/z0/kUd1AMDfKnZwCGdoma4oNgKjty4rMsV6PpTdPVRu0P0dXr
hi7ZqnbkkuewAuMZAkdtqv0ujiEiQJxg6Z/B3Jkjx3X4jT+rlRrLX9xEfLsp7FsROce89xXvdQSO
WTy4yKjazZvFxdNBq568Ve+cUUYTGauR03IgzKqlwCR7Aqeo7B7G1RmJ4cXyguyIphT7sfSe0mNK
8Nw8oe2u6F23uvoUtlwCvynb+IdkbHFeIzmZ6XT226yya37T+qUTeIUfSbZhl4coOpszeZGnV23k
z4CAlmDFPwVwaEnirqHrMhK48UEeFLEIgQ0z1N/9n3RbPjb5dN366kB2SzI1bQRnqZVzCuaPDk6h
JgY8plQmhdwue3FA250qXhzW6MVyvHwenqD3TLoDSYOGdmRX/vg81IwgO82pRU9Du8H/28pdrmWr
+cw5/an+qqTMF1l7WbXUxylSkYeCXs1EfEdXH8Fn4gXhGFifC7AveX10asDTPAYjoQpIvgVMKpXT
iLnW+iU/ply1a88mRsOgicwfo/vCe+I8RNsmOTmUdR19tG8JbxEncDOX58kqQ4cpiiFvXosbTpc8
Qe7PelyjdLzrtO2UoOv+mv/jz5x8ZwQcbHFUWfbR+VPeZldF7moBvkgcXhogCD7AoE9DHVuJDOne
i5o/2DETwM3zgn3cQITa9gS+Md+t8Q4O8uhjkJHJf9uuQ1hJxP30QBUdxvFLwCzE0VeY0ZgYxJg/
IzaLCUUBCPrWEXnzVbeBE2D4shs2Hja0HKlvk16KcubDH0rsEHkyRbfhP4o51PyPBX9FkIGLgJdq
1lxiU6r+D+6LnSJBud2Ud0tYEJOOFTCgGRGpmrB5VpilE0SwcAkrWVYWj9JH5B+PJ+WYhXyYNmjX
elfFz9aKMP/arJo2v9P+LTXDZ+Ih9ssGzeBjoNF8Eh8lkF0lYimq2Lq70zP5SE/WZlRtqGsGvcho
hn9kOaccWHKa8t+TFctFvTW1QzgGPUgKxFj22mnIyit8p9WmdRuuQWMVlFIWbmkSHwm1tpAsFLCw
tl1Q5s+NQrMaFlk3Ddm17GAUM++YU8Ho7+EjO0SVGSveQ/T3HLxhY3GntvbCQYpjfoyC04+g/kEp
WK3flu5DhylhNwVNAh2TAqO/wzgAvkiuHBDkV76sGMq4hw8aw7v/O+Y2Po/4kZtrRCqaREdJX4mz
YB697jD4mEOjnjQ2dyAM/KVxwve/l6VBF132XY2bKCjj69e/rWzrAjzxhjkSwx5VYIIbi27alvLv
JfR1O8ulgwQ/lr6GVXT18jfyyHmHCzo+K8O9CHBTJQCJ0pNE3znwOG7nqJ0a0mBh+XkHjCRoE0Jo
E1yVJc3Btf2217OG1neQqeWrD96m8cBp31gXQkR9y19oUJMFhPnS2IdGYsCjZqJUlUlvs4IovFvR
XUOHSqDAGvA6QJilQ49jAw4bEmdmVpjjtLXh2dsHrNGQPsgRP2vxCOBB6tWybG3k6w18LxXYSp9o
5YxZd9PjPCNOR2thWt8J0JZknaFPT9FUKc9Ag62Bge4zG2/2IaCtNvlrb4b13CsGLQ2TBNonOREi
6l2ADbNxJpIC40pDnLF8VKCILcr6BLwsUWCA+KlZbdYr4C+IDe67eZk8//9uxaAMOx+3MI5qLqW1
2TiY1w3y/28A62gHyv3tmA4t28ncpxlmbZ2VYO1rJsPgEzM39Q+GGOqPrdXQBFoJbSYeIuFg3qi+
fA8xURFY5xWVtDiXWmwxhatCLowz7D7fk5OI2WmIuMuSf2Jsp1sT5/NHmfbBbmH+ey8FtRDKhryH
4/3yIQ41or59NsGA0RDBTliuB29GO0oHKi8DBvpMGBbG+FPpWTht2Efds1lbL5OYutXXDzxjcq/5
tZt7C4jhQLguu313hKusdiQMg+Uyhdj+IX9mJ2Z5I0FbjU/Cd3AFbWYT50g23B3sodrHP9v6B2sA
tOHYiH84fU9FCxGp7jpnc+14TjUWcl/qbDkdKyG0O6wrdxEsNvkOEfido8npB/wXP8VRlRSq9L0L
BjGVOIOe4whVbiACg8gWY518gjafgfEgMvrokg9U2feECQ8TXU/BgVs4CqENR5hWvVfj/Nf2eOoW
HZgly7xFg1Oega5foP65DopXcuZnMmhL15oRRW0jVrcyoJXLFZw8x84K1cPaIgxTaV2zlfIJ5Y0V
6V8+myTsj6gnRntwPG7YEIVoItSeuywHl0hHXPJttAhVNGK4GPzi33wpOugjd8xP1SgvzlYRRmU8
2WPGTXWfosz4vWspw0L4RCWZrVcQFP/X5ZDqObgOg7xuMNslggjl45bxhJtKfEZo7BIqUZRZs7WN
Ne00z7w/ZxzrNa9TSDiUhwRMKbObog+uRG5CBJrxVn065+0NTDHkK0LVQxXwlJDRDekM9uVzysPi
Dv/qI2ZzyHhxJEfdgkdaP2Nyz76Zf49HSgz19HyWvi9cFP7SpMXVpZ6GnhjphMHyl+z//p+PhICG
EVwA3aADZZuAKPgVBtAAXu2NnaOM5G8pXPzIEbYgcUCbijHIc9QOD6jfNnJ/pYa0xL1UN+PeEL8r
S7N9psUSMoNhL5OBBDEF9l1w/G0E1o2MKav+qkrQ2ugocIFTT/ikViCs6nRzxIU1kx/+A4u2MPCQ
Je40R9Xj7Rr+Jw59OcHbRZ0z+IL27zfttrUOgNRAaguPkfierZ5D36sTEYwc4JGukulwn6hKpFCv
jJqMrcFcdQGXuUG8uEMpeJpkBsHjsdzx4U9fqm9bUZ0xAtpc7Kg2dE9GujCnxwHF7lLXqvZLG2Ei
Z8DLW0h2NoQQpeOelvm+Ig1NVssZsxuNu+/a6kY1s8Cb5SIVRKOUn1inXW5EETjciqTKYZLGa8oI
X8kYUJiAHfNprSL5CHNpswQJSlcdr1vSicY15tjPgF8F/rt7CR4xLXZaFKaHFcqDEZHO+Wv4FAP5
C/Bo5nvbQOc+xI58VQjmnoolYZviRpz/0qosyM7I/X/W+K8mWU9G0nplVlCbEkJJFcjju/wj/0J+
ZfOVfce1L+rKhUNaaU6EOMc4GqiAzx/ZSiDx3gqwOfs/PBGkgJ8n00B2Q5lk1hNHPTB9qgAeS5dY
OZaCMmGQKqOfOSH8GnnfpPcMdqcPHsOdn9qrsxtEImSmdKNbkCfZQEbCzd59/kaXdR6Ap2FqecFW
3W0tnMs03ujL5SjnmOBzzosRRhuDlivsZ7ERFFYQ7HI4NylhJ8mXgMQrrrmBiRskzwmfsF6riwQ8
IkyAMF8PGVL6pmHXfZkm2b2TQ7888WaM0ScOjeX2UArP2KmVJk8vj6/pDyquEn5Z8X0W58TFh9RH
A1bhfIfGZV1WhMMkydutcRBuNr7GBZI3vRCGMxyULUCO4Q1y+M55jmcJTiw/BZ3UCvg/0Hzhv2ac
VZx/36yamNUd/SbwOtR1uDDRv4++AeYfoI1K7mua3l0jrL6bynPSHkAOu9eR4EhRCNFJbUTpKwBa
McmASJ3QR2v0aOAf41d7FXr1vGGsGKou7vSce+SZ2m4DQPXlhIqV7KwHmJAxcffaNt4KlHFLYvbl
zqGSFBtWo4G4fSNL7pfChBRwKMz1PsmG0SwskGyQDYHjq6tswVew8l2VvVRBZPasdmkPSXXUeoqE
g5JmNw17KQlViuiXdTtDNRZXq10JVAnrNl6uBY3Trfl0AYh/zsgnxRksyaeh2u5eyJBRvczHXL9Z
nTqmtTwA0m4GvUINdZFc4h5wpkIaaWaJlKGXd1XdOm5SzleSbrvWPGE5YiMekHANHeSouxMTgZZp
M8x+AtpIXQzIUWMGlqAtRsxHNfogUEnGfOZSgLEOEmEYuKhBUDaGFIPYPFN4kUYOOwM37oMmMFzo
k8mjO6sZLU0ikLQ47K825VeKZJo0+oHTICXrYzadvP9lp+ixfcSg7pBRAhKEIN/GaWuujDcC/PEj
8zrLmqyEHs5OeIEQM1mH8Bep3EkemDFyj8n7+spD61RjnM5WkhzGBo8OAKnwIQDMFkrSqRmKDi58
d5M9LDhyclYtJAC5NFy4/Iw4AKfzrjJxAVsltPB/9nAO9D2LtwD1qYwp1ee1tihAgOO7DrF2XCce
cBjc+zHVTqkIdun9ISJTN9SMr10UE+ifiXQcf3v9qahty0+dFyfjuiWWzLLYWH+JzG8Ziiogr+Cd
RR38R+Xsa+ERmJ+BQdah2RY+TzR4X0l9VdkmioPVyD63pG13qgHP+qOLe42W0PT2VotaUJC4L3wE
wwurWFi6OsKPtFUvALb607fQKAIVHDbxVN5aipUSuwvvX8AM7ZCa3VSZQKajIc4PxGzVLlaklnEX
DCxWnhB46L9BnGacBuxN+BhYDyekeF2FkZ4g27k64TH728MkIX7j/2K/9/MkYXdddBs16K9lIpL1
Hh7xxeM2Sb1RexfXmTtPdwMsRzoZIOGe3XOCOKweq48AQE0BGTzQ9DI7j8NC3aciudTC/p6YcH7U
m9p6TLGmEa6L9Ty+1L7qx35nKEmzv5bbZjiRKeDpjHF6zFcc8HAhy8tznzTyn5xPssJioRmQwFn/
El3SCOWdK9nq1Y8fgBrnLR1R3QdYG/VhNCHcOvs0bGE2jahsYGVMyPMCviN/7jzEiaJoz49LvWkR
sMk7Ch5R5DGwS/PuhbsJTVEc9MHa2Qv5m5dgoC4ETGOW//YpW+lPJJxWNjklEhCvVBq1cnWyxpaB
BdoLhTNRU6dHbMl6w40UBGY0WME1SiAeUVy0CCzE3sMrrajKor1cNJBQkS1K8aG0ZWGYYMK+RZdc
D59k130DviaVyjtdD+ShczTe0XgGiyk85mG/EIt1i4HLrC8FRgKjsqHvM9s80ojAXwjFoWHfeDqz
z0bhrurr2CxRofSj/MkAEAUgd+ZWEkYDOePdJB7gAVZUPsMBHRRoJbf1uwcEsmPZ9hG0q8Sceiup
0VydMG+U8zLZWfJLwjsViLz2JZMHkvyIVVrDpXPHJSNu8YwC8IZOAKhrE3yYizV9pdxoM3OwHjiR
1/Hqkia/Kp+xLQEXuyFsC08KbW8YgG1RPckVVnEvTI3NLlqHm1c8HEu/uOJzBo6W7Wq+A/lEMx+w
zEpx0woSUM5uc5cFUSmofHnuGDw14mjw655J+cWZEUAPAS0Gs9aIeeZou4AZztnVSc1ELcc/t+B4
Ds9yZ7cdFo6TB/6O8VAB7BDjKlbxsKqrDScx7zOSyYzEz5pPrR8HzEEdkOgaDFLoOv5hKBWquERp
2GGaYvK6EEVi+zTmOldbCv/bIMd5KHZ0aSC5x67K4i3ml+2Pgzh9cHV8bdyNGfodKlieE7xf9FuS
xZMXEwmeNC3yPW01I6O337VwPV8EB52EgaUGkVWf8EZRAuU+Kp+6n4zrYYSjHNZKKxXZCQG+zkPs
sCN8O/IQh7sAs7R172lU0DWBiVFDazCp3WsD2DbeJVbP/jtfzFHHyY6lTitkViV/saVFTxdMPUPH
HbkLjUhLWWrVdggLmhIhW5Cpz4/zo+q8WbyjY2SC0u1ogzC/K4rd9/97VoKCLJDNkLg9scUUT849
fr9O1J9joIOyeHgX4So0Xjwh7QHy/HsQRscLBZlweT/IXq4mXJVrgmfkesB+sXz+fAsv4YyIOo3S
Zec/LdndekJpxKznaEaUT2hxtB49+TZUZe1a5AHzaQ9438v2sTx60hNe7N3i8yYLzN3A7OrgfSih
IOyh4W4xFnghjDF2VFt2VAWQVnjGAEB4PaLQ1+46f7gE4WUBVn1332ROpcfnCWT27rToGdaAbXLj
bE8nRmbLbo99kIfsO/f7iLKCyJ4nTlknBWz6cuR4KzjXWC5oOkJBL09Dyaj1JQSxBNzUFhw6m7Tz
9C7urP70+2AkpPWmThy6vYgqOwFhpIVn9XsYadF4VFEMYKmdIEMJf6xaLraI9+9+3zdGM+a9muc/
quQsVt4cOys23Q3dXlNFmYUMjOpLvOZS2z9E1gGiWFJJvZYeaDd7I6UOs+205rHo/onE/DBfFJpH
kQLWTiHHUIJECeRzB8MhPSMab3DV6xo6nGhERrn1GMtL/36SM1kb/KraBJ0ZqCDJl+HdqK7pvRsL
Kz3p39yLmT5+f8szCrRUGLns/lmtkY1FCMDIx4gxoXv5xHDZLAcMtygaS0XBBvaKcGLohXwz2n7B
x40/xeNaYvCRfFgHcvxpD2USn9U1UbkFDj1Tb6eCKDhOXgWhyf77SvrxEuLxWkh/RdNVcEEn6Epm
RHC8jZHTmJF9Nkb8gXmcmCprk2ufe8nti1DASAKmmlL8ZIwg8Rz8d/Ee9k+mWW/GReAZaF507fFV
q8HqkuZHur98ovb0SeEv3TsSeArtlhMZ+HkfAROWdHg1CWDVeeAbuHJa9YubeMYNgejRraCO9sl2
R2XQt8RxFKUGKh6er5MiMQy119HqYBUJCZrtnHTb8evf6ZsXXa/SKUB/bQbgjvc2cZXC9MuOOjpZ
jDfCFlpU1fjzagxMazAo16uXbyuKilQ2rxUsgiehbA1tc6UE9dR0woGetMx82ShfqDAAFbt05Q1K
RDyJqFIC3MnSrseOCBPIuWB2RpyRhDQrzYsPrMSQuXjxc88Pz9iG0bMJDQhjmGtMdPf/oWc1BJ+s
AFJJ6ueqiorue3Fk3IVh5twdQBdRG5Nx4R7tikgJflezsWxEo1L4A9DVm+kvXiQN7LtnWPpzg87E
9ucr847d1hzyZTvNtAwoFWoYMI7ZHtHrGouFlVX4+4S9S90EGKc+TYj3EaT3d7RjDWAKt404uJSw
9kolAV/EwyGtBQDBtc2OArTc25omzwUPl7qMtY+ffQCqIvenIjf/WWvXOE0sfYWlLvagI2P6qtqQ
nKRrYOn1tA38WD7WbxK82coL0RdMKalOHlWl63P94Tvxoz7z68H3SLuWUKe67HZwrGCGvwxaf7Wm
lIoM0dROn/dl2ISjg6UhqdsS+HpUKQcU2qMSje3OfRD3VYUHW4exKUE6DgstJQNywEvIPCWF0byU
6Jr+c9gm5qXvripPAN7N+kjxMag0+BBRIPXl1sF767Y99jlhIgAwXlI1J3vcHSWZxTz6ocsvhkhU
SrIPBlumTka4oRqzyhiWnI7VSY/HvZ5XXYkTfC6+gKwQwQ+EtHdFbVdH/ug/ksCbdammM8M/TwYn
eqfzGlRgWiJdiiX1zBXwSNTA/ObESFVPePvQFfc5ml2xr3dFZ1gONs2ofb4RQGfmUwXOsJE3S6IY
vJ9JZmD96I5OS+803ktbdjeqs8kuS92nRpScBdozBcje0fiPuNyTjASzeI1gSr7i+D4jdFaT7J0u
H9eLR0/zTNLqgIcWd1v5X6FVduiDSF5zDgyUH1PNfp5SnkBy/T4d+b14IBiA+sXz6vz5QFQE9gGh
KTQFMvudtqCUouV04ELZeAWW5EGcMhenlWzrdRfrpOHMi2VZkK68LvgkB57XsE2xEjyK1yOsRxCQ
ajIHMtq/ZDWf49vVE8+gDF5rr0rLWBP6gPzmxpghXkKJkAw1cF4TlMaE2Dl3h0TCcXwgggCBATm1
31eTWYF9Uh0/gYWhkDw6cLaCnmn4jo0Hr0043Z+AIJrQgI7yOw1XDXLVQHRb4aWiyELH6tMB9KpE
xIRLUT2nXBN4reZNeuHmFA9FS/XIf2bHA14YqCyDpolVeaQqengH3OioQ3PmKsDmTnEKkv6FwpZt
nyn0ROovTUeSm4j/GqngalLIrhbblNjmd3AZCEBNCwrI871RsZ/0oCm3RwwOWNfXI6xVpdg3Erlq
rcW3XitZaZDVyYTKUQ5jR9pLqOtO9VRY5ZfPwCo+OMA2fO4zDGYPC0RPrLr73bf94VK3oN+F7yB7
qW+iq4A7UCqKAeCPEq/71hIykfgjcod494NtlhPTlOX5d15Pqyxj2d0VMAtGHaJdaUvGk1BogeX/
+JxaHfFaTmq2MR/+QthwBw/XOAWKD57KpqvfU0ZJG/Ax+wZDGBX7PH91iDy63Y1avm5ZGbMDetwg
1I/L1G6sXo1IX6gn+qNB7Hnfz83boZwQT/1pgsuTMJWlWiXaTnK3ZFmfOd+z7CwziqtphHxwIv77
AKqX3zwc9xWWNRuHqcqjANXg6bd69YIcTCYJuryzhszGENlNtin/IY5l22wWvUC51FrVgU64P7DM
nDY2zdAh4hrnCcS3MDM1cYJ9Vl3RFy19IIacK+h0B+vMt5t+EpqQvBUpCQLRq/xLw8Kp3UfzZ9XV
tGJJ+Sf4TDbi7nFHuWsH/auHEVry7OpBO7YdhwB5HEK/bGo73ujPfyspn6m5668GLW9jCL78p/Me
IVZiHGBFmv5Lxb1hTwwBLGRpbvmfVkBOx+NnrdIIFMF9DC5qvYv+NHXZ/WvQwIINlGJiCMKLpxkl
j75+3nnFOpKEORtD1Ak2PFr+YovvPaENGLQEUlI0Krw1/AfQhTkpKq/5Z74Uqur/jR9+iGwhUlPe
fejSKYYxvLBNNlGOyNrXGGB/Mny1Zy0PHh/LVTNhYztW28E0RvluZW5e5HIf9YSu/MxlEVUsiShi
NAVAW13pVPKQoEbXr8NTgl93bmAJ9ilsp/56pL2Ld8FmHXjpGylmC5qeWYpIcZRzKONWhkH4EvKM
WuaJMCptzhuNtB7TFOmEgiDJt1t44E8MpC/FM4+4ayiQr4AW53aUrzax/Hi5wuMPt8QvGkgqsJx+
ltoN0qyMk8hMoJ8x0HQn0uBJJhD/8BUZNsn78V48O0Drh5zmN6lmHMyPvNCmoEmvhMQy2rqsU6d7
ba0rK9kz/PuqIvEPvR3EW3Wa8K0iRNaSHGijiK1fZPf6OU0r6Ww2letf7tpTR8al+//cNkdK0QLP
u7ribqfG0e17JG7wQD4qAAMA1VIWmaFBkhOkUor8CXEdJOG48ulC+jqGIaG8o7zz0/Y06C00yrM6
camtRmis+Dal2NFzVcfepNjfbIw3bkPCoT1f5jKW1qTqopSPAjlGUuUoPSKPjyBq418lBOrUSE78
qm+oMO8L4m0krGBKjI21bEW1A7G9E/uyzLySbSxMXfpPucVOUnmdyt/uj6mgkFdLeogHH2TCi0Fq
ZCyg03iEVb43PSF1YchANcHh7KQBiCxvGJIF9C64z1PUselj1+u8KsIuP0VfRyVxQGgCOIidTanz
59Ytzh46LLdExdw1HPtQOx0jdJR6g1Rv57hptkLS7wi9t0k5w8rgOpjD7s+IWK90Rtgp6iJX7fuk
aylvh6nL21Sk43eaImb2d23tjt+etpJ5HlWlyv96fgj+LO66W7D1SxSFge4/H9ePuBonNH13ULRo
0HAxI5aQZaWENA8hajjghDEGnEkfYZcoOwUHxsU4i5B9dzfks+F8AmRoF/pCmHYIsIu4BI2AAPv3
1ih2w04rkQBJQbBvjTuM03Em9VI76xruJPKXJvdlcAwpKQGh+h7ajZPMAQgJsgY0KBTtDg6UFXWc
LNihKxze/ZCF55NJvJTWJoNYEITN9oAzkJmtgkcLrPoWEwX0UiO8kMmDAYOsOtmagrwjYH5kP6Od
UbCoFS3IDzmRRl84WydJAWfKpp/baG/ArpYVXcZvYOyTX3SBype2PzbXgi8PIsY+hvaVqEk5h5qi
sNdGIYV5ZJvoSm+n+60GoOVMNIoQmMfwRQM+w0amVJzsSyM0CBALxBtj4nA0ArbY4eVIy3IxpqSd
+i+h93m1y7kiHsMwhp45Cr0LqbzEDf8UUU2j+2zVle684W6wxX3NiDEbGT6u/4ODsLXRTrRidOdU
ppqUcPVnSFq7ezxo+6nLPXkPspfZrl7rxFXk2IRDG95M4j4JCs8VfW9/vxdyqpbIAk+1BT9U43o3
XNWW+Y8e3Kgec7XIAACavQonHkyv0ZGP+gcGhuWAHJ2KFbNnv74rZYNiVcz38YhBzqMlvvb7NhyM
MyJLLbuQ9uqPibAY70a1MR42oCEJuZ5X1613F3j247p+CvybmmWvD/skgJqF/PheOhAmM3sMtruG
OsKmSoNA8r1TD+kZbGgknqxu17PXa05iQvQpXopDG+g17ACcyo/XUT4jg7xE14VzX1M0ro94CaYN
kedSYvqlUVYlTlfsVZGCQFa7mF1xFzAGYKFhsUXp1MWyN3krauHVvYZHE25hipxncGljRxDpcxWk
r/JVtU2pCxnNGwg+LjyBiSwauH9eEREw6f2TVRi10voS+NwvMySsQ7CaaJwAysvkPK8gqJjBk2sc
qz3nArNdWeNZCXUhXPv7GlPUGrAGp3d4Pm7QdIG/C/LO2h0eqnoH26XbhU6+BEZmlhyaydxm9zlD
HBzZM8HJfsEiMTFFGVhp1AEeQprR04/3EJU41jx/jSWgqBIW1+dI9rIhplWyVpHv8s2kU7vplegg
KezYbawfo9OeuhOIJ4eIB/JZ6cOAqFP39jhZG4nIIDa8EInuMqtTWWcCU9Vqp2Z7uo8blFhGulP5
eHuX7zQpCfTq9RYNSG8x1tmaygVFmlEppmdOUFEoly2wiqde/5jXQxTnqak2z0kJUy8zi/lOQKup
3p6Pn1kDODQugC+EFZMhqve+EXtWpcAU48x7EsMu8CywywQPchxGGqBGaC9F+RSwR9FCWDJuaZ3A
JAejXmoKu6XqGa/mUuCzX1vTME3ETvyKx0BCwkcw2AUhHgc2eNfEM4MrrIFvN6sH9GFTplRAF7YT
KH92V9zn3Qc3V6aP2076k5nty6MB4zCZtNQm4N/JZXvT9m2IdqYEy+kaOw81f9kGyISJ1VR4Jb3c
e/dpWezYtjSQRdDWVheaCpCUyIoVE6yTMpzfswh2KVcbOSX2BzY3qgmNYVBQLURzzsYj5qsZ0gyB
d1/PbMLyURZh+HCuglCeJx9cggcFg+c7d5zT9piyDzRpUdSzD+mpAbSVzsaALPXE8jIyijoRFC3n
MiHAiLEF2/MWVAINjmUAaj05sDKbuBBt80vcjOffhBbvoNueDmUONr/psF2aTnLw/Xe3F3SHhHy2
sC4DbYGIWTxZmnxlR4SjCqYt9L0y2A6rDKmVtat372bR0yFwSwKxKoqPIRBRpflfoL7mCmCGCIQh
Ai+5H9yC9H2uuqzwfMllKQ3+7IZKoBuG8phU1CAU246SMaYjUzdTzqOrZkXxzi9WYfA9bKKMhwn5
We4Mn5fFXoHTfYJUxk7piGl5DtX9uH5p28ErK4tYToYzadfDhNlq5tl9tIsIebypriYX5igQ03E3
dkxrNDePCVjLwAQnDCNwvj7F7w0I2CZSfjXRJfObdZfEEqbaNZ4fo0LCI34FyzQLJouzh+QRYpqX
UhK4jz5reEdkBUzSfAzG2n1hdB+hUWpCzEX+4SLP/OXb+GNrFaa4Cs9izKelIx81Ba4lN/qkedqk
SLB5JQNJ15Xk5lscXtjRAJm6Nmm0m8b9YLDhBw+0gZX0ONIfmWAMn344Lj0lryxCSVzXuaPJ01I0
o1elN7D2PO1SM4fmLpIuF/5yP++IOXdUZ27J7Hd7+Fw7IsrGCXKEtz78HU/R3I6NA/dflBXV+KH3
WRv5CWpFophwVF3T88U6MXO4TZs5/4FjGYsIyn15fw2BXhLj3IoTQYd5/6dY9cmu28Km7Kc29t2d
3yzuW0jwk8Jaxm+w6xyEIhcbxrgHZEcGv7f8la1uzxFVJ57Tn/8GkYXzhsrkazG4jV0fHrw5EaL5
qxNNgDHf0CdlBpcsY2WKhOxqSatWXWNYQ+gmglo7ffTawEscNJwGr2hvzPEinrV65VwcGwq3HLw9
3vRZcNtaYDJpyXMRBlqgvclvWkdfaFeHjFiJ/vAwG24T8VAjMJuvem5nsJupdR8OnMIIferPnvO3
6KT2psK2QrnRyIwhvQJugyq9mpPOnjquZW/mZhQEf+Go+jplzoGoflA7GiOEuK9Hc42Q9UpEbaZV
Dq5A6lOFGCaancjQJgolOUlqS+LeU/vsSEuyqTwG09Zo3tuMbjQmlmW18jYt/3yyE1wbt4E5ufnk
xIsGTlpvYo6GbxnIzgOanA2DfV+MxXGQReN7RgVx8HPI1esn/a6y7NoLzQYii0W+c2Wif5GDFe3J
kptlJKcwtIcdVQKJ87Pg9+ljBmuNCHe4HAUwWL2IqGqnoLR1yFv954mfQAkAtaAvyUI9aPijI5PX
uGF3jECzI3q+z+hbujWqQXnTMgbJ1m974jBEzSbZ3Fof2Bpa8C7RmojDVVBQkKumn8yIRt6IkJ0O
/t1S2KJy5TcEW7vBy+kpFAjd5MFiD3FSeQJuVLyWH+1mky2e75kJClqhQtLCF5r7qoPkGfHtazHe
UDH6BrBaOdcnGCndMG+lmCGqRF5/WFswjUkfyh5x/Y1C1BHP+pAdEZ1YyHXpeQNLmcFborwsqOlY
KRvtG7HGhj+lolPP3X5bMTYyoGArG8T4Vyb5/6DfTqkcRXTEFGggejmPAh11n+Esn3Je6cKDO/PG
A9MCkc79JSSxxYzAF4leA6WwSJ6qoVxlNv+9pFd+YjO5FwNTodjsIBZjApOdxVRHSkqUzi0mJ06S
AKHdtSf8/nWW+NYw3d1pKSNAPE0V/X02fw9/l3YpSvmbEhuOPocVDE+kEmmjHdA5n4iBYLjS3XhJ
cJLCq4LYaoIp2YO9dLNqDiuuLjxiT6Qv2da6wGw5/D4DpjL7QeXiGn6K6/Z72fgyAf4ZxPocGyeq
OXzuzHt3FUsP4xYG+lzL7dDTuOcKtU0MygCwwMN8/uCo9o4TI28fJXY/uauyuxK+xLp1VZ5PxRQI
rdjNP9KhrcKrbHlg4tertQNYTtMmQlyLP566gnd0zNpP47tvlMo8Yhre7b8xb9Pre5ifiECcN/BL
XgeqJNll1SIz++l20LfNXuNGcUzBEWFsVCqVg9YaY3Bn1Juf/GdX9/f95HVSuniFpHcL3LHqmoQ7
B9WzHVAi9jo8zJK494SrPBR+AXFXwbfR3XNRyEVXsLTR++WCku/utbBetD4+6GfwJ0yVusD+/SXY
+/Bkb81IQ2yWbuuCe//hGhOnE4T4FDdEXOx0bTHjba/ueg/VL6tBWMndy3o5Ywognd9jQhWINF0y
Iw7DPIN4ang1DA7AgPOn3mvvxY3RcJ86xUWTqC3hepwZ455MSHnuieA+t9SF78sUlqxAGgZBsCp+
ni4LIcbvhQhs4Al1iZubALzZsOYeArDas6M6/MNYu3wn3o39Xqj2bX/WSdjCef2A7SEVlt8ZYugg
NghYukyArBNRrQi56eK2mYqMDRLx4P31XuNW6y/k4aQTYq4AHbXQs4O7RhN1v4PSR8/XpC5WkPsF
I0tAu3SSRlcS82mN6I/p9jOSYFhWwdeu15zEvFO6lB8r8ly5FI8aJp6cvyoX+w7hb9o6FbBh12nN
ItK1OtHHE9C5RkGUcztJFlgHlyCAE0yo4tBgCb7PQYSMKu1fLOD6kc4Yj4mIbxF5u6IcuxZmJE19
uBGq0S3CrEtoqskWUrauu2pgYbXvo2rjchEObwhZLgUjuaG0ZRnkKOeyp3PumyZ4PeCN31UHFECD
AgR74PJ6T6iSocN+LrDQ1YSNIjcPNfCRKDz8levXvGUBmeYyyTeYm/0U3jZwuQmsT8PoMrigODsJ
FeKvTmuNkJzyLWV71uoK9zI1QACNg0tahjY6WnrOSPIE9DhJl+rQTi4C4aeaiavmQcRa6OcMFc9F
Ed9IyeqtTgO+OG3MvJfxJn1by9BEYpvAOvn/9lkG2DfkFsKthxCQdB55XBjx4kW7xehyrFIyxJ1/
eA4ATgmEYNIoIIW4um7xhWwuyqdWea5/geuYNK8ZV7n943rqSLa3SDXEdbFzWULXTvpZCBfKdJT5
miyf1pOnK1ScelkwwvrVnZM0oJywymr9MreOgjbryBRqQoerKsFnHWhF/RN4SGb6Ymebtzo8iyiA
qAxsq2DnFPXQTIauZx85qIsNSo18NZAPRPJayKH/Rfc6SaglXfaOsDruY0fWxykbfhpRj58sIJ7i
DMm8alQQkL8KUUGNDufpS+FQ1b2wEWAHos1ilmT3JU0SOWkceRu4AIcNkeyyaV+0NRW4Ab3R4ejP
8TNKmfRykdys8TRTgw0+1vvPMBdkoah+d48ZBojpwMtlV7EIHpKts81RMdeJx3VdsM4qI0ifRXQT
IY8pYndIU1WXUPrC8H3Au6H+BP0Ewy1X39Fn2d+bxuGOT/35ZJSLxtBkdAgEVVCIGKqMTE2cBcNI
UOfSUClvTXsB5TiuZRLCLixpbMGGz2V3Oc90Q+eS1rGAgDhZfcgVejabyA6CraWKrjSbVHlCx0U1
j5qzfRtfC+jhrNQe9BOdKt6CLjN6Ygn4dPAdmlQNGQfoPK1CNZUUuc0Z0Q75FRUvcFpN8b47RyLF
URQYWFSSCrEX0Nt/iJxtUe6TMCJoe3s4FeKxzAT6tTZqM6axGIVHzl99NVq4LJTaHm6TczRAyjtA
+UaIficvHH5ZxE3df9gaVj3ErzOP1twOvs48lckpb1oUdvuRrR37DB3UsahXpFYOba2OQHHe+26/
1SewqCTmI/V3i8dPNEgfwSZ+NN+YgxdwPCgh8Dk3zhjDGDVFBXD81jtBSW0B3fTWPnSLzCe6YjlD
wa3PdMQ99yLSG4LiAP2g1s4e6y6D71IjfL/CKyih3JhM6tr/GoJiJx3N1TF/T25vHsIPI6o4T7Ht
FZXytVNaV/DTXah5uQUoaQePPb65/8syjn8UqJQe0VXS85onsKJiLBWqsHkH6VEjGLdVpQjxiGrO
p23zhdhYrntWHm6QLJxe5Fytmi8M0hXBUqDukEhitVwj+5JKX6Evic1QDRhc5nf1D1VEceUnQEUd
Kqx/CTS1Bhdk2iOk5BCSTIXDUYydi+65dk1PdgbpgQW//Pydpl7G1iRCHTQ7g5nyGzfJKd5CSXcY
mWHprjdLQxLCpMdzGGKJ/cOBgprFrvSPsqy9bm88bGiHjVgcHed2xeJRROsjQlFt+jo7JuMcQ7xm
MjepU8co8WkjsT5FleyE74i5ta+QY03g03ah3GL1txCds8b3aMX3YafyZrRM+m95KyoBuBtRpL0o
523U4g27pZFlMBQLHAglur44KupOodABW6HMuA7Uhopb+b5PUx07gvApfkBTK6NJFVinNvAEVOFX
YfnHancVYU22fTxB4/m/9lX6NEIY9bl4cMfI4yFxRxRIEEBC+X/j6H/vGe6QZYAsiGUXMCQZ4PBV
gHEfvmt2TZUaDsVAtZtrexRwdeZhcjU0Ls1fZlSaq7GOaUrBW2TynJWkDYMysT5nOryW5tlHxFC1
894HQwHFZNj/eLGAPwLqAzHrdtIA/yRpyDYTU7jSwggsqB7mYe7i7WnTm76nYTU8pZ+TiO1JXaHb
PIbVYpAytE1iVJGiYfN/V/WCFROvdny0aa+uyUDLQzX/o62GETIOSjRQ+DVZEppQXWrDFx3SQhk8
T0TpKbAOjvFIipuOhNZIZPnqxKswFB9l+tSfFO3+jM96uBPslPfpip0W7+zKctSAfnuPx8Rn1M5T
MeLfHSRShfVSlzNSZ5O5yCFUsZDt8ff4p8ES0y6KKAnTJ29xvNWO3R+c0LJsPVFxHPsaNPC+Lnto
92jRqBaOZ2J+PU9nGT7znqndE5P1RZT9URTB9xGyL3A944REMzU/Do+Im3VjozNfsp+2DIsO+A2r
SOrKqA1u9a3moiS48N560NZzaiUHqan4T2apeTvvB2oo7Qx+sUcFQKsY7Yqf/dioVl4Wk5Okasav
AQjjxkrx+9nvjKKnQdH3c867zoFn8tmMwwCOj01CWRINJQ+l5IQA2uw5eORNq4/f4D8P6yR7XQPD
UD8c41CRP78iK9HXsgkrteL5GFsXIbZL82YvqeUL6JIoGquPsZnVhMTTpU03aOHrAg14Un6NfWCO
vcsV5Y9LMrh4U6OiR5xCdX4sjrPE7COlESutfnaJwt9ce3Xs36sTUN2oqvilCm8xfZWKzGv0qVC9
MV8zXlgcrQ/1DsFGxi6M43ZPogShPZY1cxRWCi4d0hmbIvO6mhgQpvPEEsxL3AhLdlxzDENTL1ce
X3CVqV+xGozyytTzVL8EfCbJEpNwtUuAv8cqIWWSwSFAMTQlMk+aG3jro4Ab9JZHeyHgD1dyibnn
lKAEPkptGjDiPxinDrenYnGMyFlUM/3sV/uaEuVIi2ReIURUd0Vu4zfKp3Cm0OJ+aJ7PPIv9E6Dm
l8k6FT0NlDqzNaHexZX6IPOSzT03LDQtwhEOcfE2Cwv+/awWJykDVX2KkJQOblR+CALSlaly+05b
J/aIzNr+RvlEO8opR6DFwagd/L5nekHYkDzPvZsGweLQHzRjxrbvDzS9X+c1OoxmFi+MlP8vrYZx
7ntF7QbCJ5ExTcxXtfKk1mR/JU/3isW3B/evQujt/K1dxjYnbsZabBmyr3cHRV4krttz91cTei5s
PYMX1y8j0/hPXd3hs10Pfv99yKxCfoxcKxD+tXaN4MjGTR7PNx9Rf6jy7rbDj0cnzGQt+Bcar30I
rC3mnQdF6KLQNETLV0OhKOkZJauPRHeCqe34RxStANjMoMw+TQp9e5tHASzIjnKNz3QthMQhc5bE
RFHGGcmmEqXLORcCw+dPnIjdsZW0PCpw8UXtrBA5p3gwR70/Q8eTKdi84JVOWAdSOoEhBQq8FeSG
mFDlujAYCzQ6Cwpo9wl4EMiXbqHaSUPYXR/V/nTObnu7IWNTTvz7yT4xU7lf1uJYuIGnxQJ56Xe/
x8NY5OcnUyq4yJeWWRnaKK4oQ4/QzX4jLwFJGsFlNw06zoNgMvJBigEyxBDmr1gdvtRxOie39b4l
yptaEL35XLWCYhJb6DDBexxNdWqz3QR9OqH5AGVTjeoq/2wpXvBCnTmvzGwccPnu3EGZrP84oFU7
OSQOUPdZu260H2tNvwYbk63SSQMBgaKSDUIjT9L6xzlwI8qolblov2Zvu/vo1I3M7W0H6RdbLRpi
xMMwVVqlbdw0viqnDuexOabrgU5GbrM3Df6GPm1xYYoB6IqhBL3iF/9vNSwsN08JiaFDvYCW9N6F
eBb8jDv9vgua73WXN0ORcZFs8o+9vlxkpSPc++W6QKLn2pkS4ojfCDhC5p/sBCgEes/Un2tfrXF8
DiPjBCBt8/oTdKA+o2jiR/UW9RtPfZ4CeLnQIuyut86yd7BJAgxyRwaOw2VhY8f7V41TfwiGX6Pa
EX7OmPz5kpfdNn/I/ydqEy0ZyqUXBw9RcXhAGiXWYEaw3CS6aHssIP4eneHkjoDvdsBC+/LC7LfP
0lC7C5x9tGnNY3FhzKwHjuiGuGwI0rSbipenyKyUT8j/0Xrli7nHQ8UihasYKyzKBecREqnwxSo2
hIJFnPghgC1dZgxb8B8d3zpMV7YsBCG2MwIuDxvKFC4Ex5oSat9KYqIph0bY7tqzkQ/4f2GmEblF
Q+UGTDS415r2rqlYM61IoMj8dKvHtt1H/CnUz5gzZkOsbAcMGNkNjXolCKEKEuJvcDc0f7QMsvhG
amP0JTiKJ0jIx+FL8dyMxM6v9lvHcRnrw/5H9/GH6XVUHy/RE5H8Pv4gdgbnQr/xzgvSy2emQMYi
73ZffsDZMqFSuS/6v0oHP4Js9V8ZTz129Ms1uQpsnQSwkO0NZy/JipcPiUwBa7Fo6Xdqy3vA0v/8
ljxDOwn33uKzkWVaHVxQH4LGoxKRcJb4JeDAsdvjknNd346ZdKJunNThtxaMZX5+GbRKkWfQGul8
nU3yKb4595W/Z3K6aWr0pp4gZmrVV9yxD8RWMZmgeLrjLT+ufw0HyoZ2G/pYVwNFnOXo4M9RO+Ms
w2TxZ4hiy0DP18qsLsSGdMN+w5z669b74HkQIPHRUI+HlhRsesLoLdjdJPDiAs6R3WHgYsDQtx0K
3YAKJMVWTGSNYrHxG2U7G4fYpy5i+7MD9CqJxUFJ+MPun+J+jacOYEfUA+sd7WbAmBcJ0dtAXG0W
y/hlTyIo+U4a/5NSgQdl20NXwudldnz2ud6JBXcttoFGsv2lz2bYS+zjft1oTE053NG0i+l15lAb
p6OPZMgh+h7ADaLJ5hIjanivZEpNwEKo6K9Qgvbi9kTw6xrGbKZpHemf+ljYkLew8RgLdJc6F9if
TFGw8ez3tCS1vW3drYE6Yqv0idmL0XQguPsxhxsnEfXoz99gfyo8xjNAK5rV0TN5SAe6I/NFeWVB
O1p751pjtrnhGYYS85d0sJQLKq7yK63UTXNIo1fKxk5ja3u3bdr6G/uv5Io3pq82/GTG8hq7eC1e
tQrxTRyO4JAFgxEyFerioMvevDK/CNzkQUdQc4RwBtJ8JFFlZpEYijuHKW5edKsTpjQ3WKtjbYYM
t34bcdeevH6t0lF7e++ftKiPA1kUtLxCfJ5VHXBZ3s9ZDUx/BCcWLaAH9WY7tzd0Eg5NNRkdzGRa
iHKja4SZJiXlcIarzSPpUBFkZlOXe0Ec012KNl4cOMZNz/IREKXUlPzXUcHY5hj2waPOnq2mJvnV
9fWQhErHwL/njIC8Dwve+CegemU57hpISUnbLrvfE4uNJlJFazSvDeKK6k8g4S/4qPOR+GpNRPqt
+nEJ77xtm4xlO/RGLeKS+QA8GcJaltL8bwF6pAJinmNr00w5c4yVVjzjZHozb3qc5Lu94yonpkJ9
qe9LIzJYeGYlp/iOKJ2OK2GHEtpAVEhuv4cLq9lwp+5dGd1Pt9LbWxtK/cXzq+A/ZH3YVKBFpknN
2//cRUQBG9rRhV020xjzks5/oUOa0/KnbWPzAHzRHEsfkWvrPJps1t4xcwhXR1KKhU7nUrjG6sIp
deitlCWTKkhhatWJIt8hD72vWK55baPhEXHqcFqAGDf1+e10hIPwsmFIc5xLZRBdn+lKJvfn/hMo
usoZWbnVmlU7+ZEKkOiQexSl9eXyDJlDm4cJqFQBadXk7bBJ93Rp8j2y5OC2Tzt4qO55Rmuxxb+A
xS/AJBMy1vnoQWZxWeqCGz8xrnKt/cBKKrdYwNxBluPRvr4E7ZsC9qjNYXhg9jHBOxVuZF2wSU+Y
y76D1ehw9yNJg+nna/fqCViZHZ96cPvq2V1BY6fwCRU8JExFwirqUeJbEu0qGCzkJFU4CF8jiKNP
dZTwB3aO4cgdk+5ZzFKGd9Hem/QBQIsZ7Anwuuk3JP+9TY0QE2VwcUdN3yyDww2V1BSXqdQY/4K5
YnyUOBFgPjAsY+HtkllxWBpKuV6in7npfpX9RSIj89fZMY89DCpmpw6S9GiUYUK5qK5Y+UYJ8gdR
ZP/yxk0l+/VKrR+GGO+hxaUgCdca0YLkFMUiDlQyCUdzTgtF5fiwQQPen3kYIDag/7SNTUkVyJJZ
5FwkmWgG1aYig3ErOC1CyBkkvFXxs2MMbiqS3mQavhubmfzPmNYWbaOMcMiD/JgXDI1seeQid+Pi
GwfyDeVHUK68/wD3LGjB3B4oD9+MlPxh6C82p56AaiaH89+iM8qZIwaZfhC/gJH/MDIimDQE1dzi
YNSGpLb5nv2dYCzZM8Ifw+swUcx/UZLbgnr0EzYCTZRyp0oIS5Mp4AK+l7QMjvXT5UsqI5J2E3xJ
OmFZMNvPv9IP83Nu9PXROu8NrJToMJhgY/K+b6YxKmRWCfsvG06qWAK/UdpKed5J1e7V4KqSypt+
/BeY4aCjx2zQv2lI0LTDKNsnmKG1+FAAWrRqLc4W4p9jUtRUWPmqSgLWRX61zdSDf8RJtMJyYdb8
wOflUnRXRpLB04cWug/S5udSwG9iSisj+/Z33wl/MhKn6sMj/J4DmqJVuPj0uQn8QWDjcaDGllyD
nD+mhe6DyGGFVwdm99H2fdpZ7CYjTGh4H2OVnr72m+4drS58W9xKaqzrGGxKoK3wF1gN4xTzJJXS
7Ht5x6ZJF5ONKt3A5VDoVy0ItKzvUYcA5rgAFHu020NRIqL76GxLDJYWVNI9OzjRddxeToSoQBUX
u2JSZaHvfOYrs2GbtPTXUvD4g0wvdd2Ripr/SCzjL75plTPKYiG2//rOzQVjNzACDh8rMPr8KA6y
5pBSblb8MstYpYgagjiT4bnrrX3MZbppzCwmlxrdxhxpN5Cx/wkJ3JNGdBMk6rUOcFnPKxfs/5fW
qbTiGeBWhrua2P7ZQ8dR56rjX5JNKxe3bkv5iGjPlkv5fo94fmr5J0rrcronj3ZAPurhonQjCQbt
488phfbvgJKB7bFS01HfCRGmdqtJ1TJJjeA8DNcJQuc0/gVphI7B2/nz4xJECZA0jF7XEawJGWJD
8w9yIhPilm/CqAJNRBPcwMsz3xWe/Z+1RCJWlxcWepa2aElfcI0z9WXVpYf4MpA5uPplATliCCjN
7tYOlauLoaKngw+sUUjjLtFmvQ98kV4a7akY+G8GnCeeNPs+ChKbQWeYLuPT0BmTFRA+/XcdI2BH
end40F5YN/haRhFEZiI9J24cXt7xK6BmmSBQ9vk6IHJY6/t6XvGL4v+wMutC2AmmrjHzYV89vKV7
uJeFOfLgESPpFnEzFbao87DiY9D+zQEOJKMpLvStZyTm8N7Ax5sBbAY67D9GkMRwn7VsltcHju4j
zf7l3uY0L6UVJuMrd36QgRBQwCKMkom6bJnF/SEwPZt7MfUZ81j1f/TM/wnFg7qTmRz4kE7Fyeuc
DS3FKIYvj9Sd3HChZVOSMiAnBay1vmUkNPonG78YEd4z7YzXcEknC1huDVx84bay5s93DNTMnMKi
RXWo7lLydIQZ6c33FGhbiSTulQiZ09bnaUIRcChB4eBaDCD02m3hu5iyuKhWpmtMTxeRTS4pCO15
AKlEsoX3AuBTP6XQqagZYmCUqx27nesDMN2sugHBzcCG1bR5uI3Gj9jSvZr9jN81qETF8EIIK/ms
moY8JpmFd6Jm6ZUPb37BMxRjxs0dli+zG59x7B7Squg4gaV23T0+mFXwZ96zEp/8yQfql4PVyozW
7fZ8730FUp1XkuRRHUodFO8UM+b1KQozywOPUtl3ZsrdhgCFVUAaQqe/G9yr5KCtbBVbwOhQkIww
jrdtVl0Jg8ErE6sObfBzI1ZlC4Dxha40RPCUC3woaDl1f5s1zyUc120UhXdRpCs1QmutO4C5UX+2
eErlhDx/d5U1A/sy75S1ckn616Zwgbx9LmEW980706re9A/ZZWpzEhz2M3WUK85ZOk7NRRZWQ7sy
sMGMG/96KLUpMawMGV3bxUNPIgp+u/1A7W2lBCm45AgiuPezJ3ncu2lltbxZDvl+XRxW21aUThis
Wlra5ryDjW6Q8vQ5KRnT9HpJSf8SeskJ4ByCD5FNq6MEi7mhntZ+lqEVQgNB5Y21+oheqCYwzq6F
lWEEOBwNQoMraKGUocQdY/KcicskWmNVQtsM8Rv15rwdRQXOo5UFkhtdoECFaU9Esl1f7ObV2jKf
0xqxr6pnjxPsUafgxWC1xF6XzeiezxYHwHzZpaQMZLKgxjtgDLi6uuf7HcJN1tBKVNxBtZNIPQJ+
NxuilGcYvKkIevcK9PxwJ0KOTmM7Uq8szo5izSCHKUJ+oyRcBZAfLGP5HfZH1jauZ4fqNlRDzv55
v4E1KzdmHtyu9WbPcP4bluvBobgzQWKNjF70HgC7vJv86gPEPeuZc+RN+qfKYdDP7MA0pmfesRQl
0MXpuykLRCNfXZipgZxAb3QqxnZQEznOgqwgRyfMhz001eiarODyIuMBfajCE/4do9s5AqjUmI2C
JFbYEZwH4m2DnGg0LuoDEf5K9uVhX7RgryxXsOIwL92gBUgxysTtJ/7dmq87M9T3ZFzWqml7fCzn
ndmtlPkb2r6wT25PhFMKQlmwC05w6+YzM2o18lL8SGMH+qoJqaQVYa89Id4bZ46L72+sNsk2iMDz
b3FEJuFKZK88BtUJtBkNU/oB4WxQKMCM/KC3n2NgejkmmhnOTlJFOIz6yr2MHum60Xde80U2YtM7
d6/0cGq5ZhoqMm+pbAwjgr5751RgJQJ7GchH7Bfmg8cOB0xqM3VHTd+lCu3QW7+FUW2ur75+6Ypt
zFaitR/Iue1clSCZFip3PcOyAjFWQR/CMpnLfOz0PF3mhzSJozJXSHkK5ZHRAa3HGkx6zHawlk/O
0NyBeiGlzLJ3JdbWjG0bxcjnINpWfTBJrgmmMjQdvlSen7nEn2jtu/0X9vF3B5ZlM9dRJq0QVa3q
5/6cUujyw9KXtL/G8J90eVwW9OZI+/Fs2ZLXjZnjjoGsGPZiCevgFDnvSmRSv7si5hjxPxB4JUXr
P2TVAck6xiYP0j0yTgOYycohRqg517EDtsSxhpxNIyVstaPiorc16lA692OcquhsvO+GpMJ6itxD
WLTNXj/OgOrkj9Vu97XjX30jisQ55/rhLyvXLPn+pMx1WARpvGAxnGff4rbuKEVhaKBLxvB1cLOI
L87HP/uwjLJerH9a3/hap3u0jgXxhD2RgyhLunZbrNK5c68kRbVYfu2dbQNJOiousPJrt0Ap4ouZ
VV3ChOMJ+qypYa/gbkNGiY7UmRwcD/y5YPtsLAauM3voUbMNSZrCcyAY8Ldp0CrMu1hYYUlkDtYN
+GDo4Zgc/Q/pUYv4+RSHlp62+UeJC+IqSaQKTvktBp2hXRyGE2vJXNZYjd4Uz0Y8ZJPMpAOXTsCf
pRTv+PYFoKCsS+++1UbT9iATkkgmJ/zTC9POAgd9BXDnVRiE283ZH7e4ejqD1L25VymDd8s+BAIL
wkLD3cHDEcfpeTIy71L+Jslf5+lBW4fZVBCzk2E9Jbez+AIf8ZjfX1sJ6j+sD57iqXKPn4yGrHNk
pI8Hekek2KHjJW0nX4TDSBtlgGrw/RmHikq2MRTKRZ5eghxOJfnK3zLXww1Kezcn3sYdjo5bnrDt
Xaki1iJEhGq0rrznQPproS9HnbE2TqBUP1vIoUbDToV7hp/c/66uK2VfwduosrMvl44pJ8zaxwc+
+JfDzBRIz6yE8sg6d+Ll1+7SGxnRe6UTlu4EFN8XUROCxZVAg4YQExFk6y0tkCWakIh0K7Yzmw32
SrNzIVSWC0qczfGQjGe8qHVmZ39rYRhz6VO5GaI1uPyWLB6TNAijzVd7sJyG/pwmn4JYiu8pI+Os
MORxAd3M3V91BOvXhjVwKwwaWSmeH0xJpSHKTkmvTc92w9CnWfm3L3GxmQGMrTBKDZQU23sjkV2W
4JRLa1mTkc5bQy5Dv+WF0xWKDhv4H8YlqAq8owsfy2NwjhRe0V7orC+ZKWrjVp7O/M9J/Dd4YOdd
YdebRMxTb02+lUk+XFiDOf53jLx1EY4AEQSOCjwp4/sfdxfAte0LWl/JdHC+LWpZkVcBRQA2ALqW
9gxk1ATXriHnJJEcsr8tbI3hR9z+wnvWIgObTZ4t2WhdzG7XnmYBulXYRYYNjxOxI36AF0KH1zEL
cZuYdPM3oh6pP5KMdblUbKo1Gkcck2wpopXkfbs7ZWSnL0kzRhTOWSQQehBd8MV8tT5lYMZbZeiI
z9twySo0difCPAe9mM/bdoHPOfty+MB+1LV0uDoIumFbBhyIIP6h/q2+rC/eccTx0vdZ/h/kzj8C
9hr2n6Snm16QfIQqVu9G5YpTRSOICWxFISfQcOxlIBHN7G7Q6nkIAa7HJFCUiaK2Lyw1Z05U1cq6
CZJ9Djnkdph9O3Z6VDBEc42nd57BeKWCYkofGz87CUTvn4wnpu1Z3N6Rp12VJkrWSH/V4J7Ln7+o
Qh1Tv7Gzdu4VN6I+kMji9BdARPRcC4qyLABm+aEb3kytqo6fNw+TmcgUnBTDSK8/+iSzqcGyUoIZ
9oImxT1ZzmuF9Gj1AxWfqogvXZYjo63vMeMOGgdd0xBqQbL/QFRZQYWMno5fqBdLe4ZakdaeV3kz
dOVroMuzWfOLtKOiJhyJbg6zapRjcT3pflN/DZeUumxET3VRm0e5wyiqkaupW5OZM8QUzgpLo/kd
/bFP+V7PBIeWD2Oc8+E5xQvuDW8ICy+zq2lG08+pRLNgzKnMXQ9XC7WrlNmSDYZfEWyUAfhdoCK0
xfdSvYM5EgQbhUC8093QyqMffm3+QKrZkTZy1lmEFZiibUjFMyJvHw83EWPV+nuab7zsI5oA74EF
8/lzFq52xn6H9pb+S0G18xDC+dZZ7KoyGz7ETA5kxJebpcz3j7ykuk35eh4xVwsdEM/Og272d+Xp
SzV9p10Dbvwnbi/As4qenU7PiAty4F3n7Qg730c/hJZ8bO3rBsgG3++SKFSog6R+oyqjdkh4PaRm
6GeCnFxgLSlij+QK2q1nZyJ4WN+uKczYL8LJ+HUMbIPsicHgn8ZBd2wXyWSQi9GSOig+SkC1Vbm0
R+6sc46bmybdzQyoRYSzpwH9cZPstUJvqRfM532qZI3/FnQ+AyaUZJUA9KNclHG+yaGJsfpp2OjM
Eg6Y5sTD2KCXz59R0Vx4KCrkcM5eNziNTcbYacoH3upIa4gamuG1389x7AyaV4FvDqrIPQS8PcTh
qtvpjhuG5IJrkTDpUGBD56AsdOxZsN2Ev83UykP6fqUwLwxKDDIgvFW3gmTWWJPIgaaj4E6OW9wz
zXcsV+v9ka0w9ZT7lvAaDqG1w2eca8RoUYfvKbeydGYmN49M2WC4cccZs0HFh50NZuxKajuis7NC
AO8xICyVMLM+3B6dyqQb6YSEVcOpohsz6hMogC8QAI80o/383gllq3nWxAr1kA+xST1jTe2oSdcP
IYNduNeJeZCeSeV6Y1UkQlmOnYJ3wvVBCkmczwK6f4ZSKrRaQWTov+CNQK/K5VFKNbEoktND9Plo
i8JcVb1mWH11FHcuF9us4t0OMD4jgk6rQzthh9oLn+r0HCogA6fLRMnyCh4/zoQDMWr/XrpjbtBn
++PavdQBxKErZvPKyxgnWxjMEY3AHbOAv6kDbcwQ6vmRloGglS/q/YMmhH2lTnRiWMyHBmycWUMc
uA4NKEz3bkVfMsxaIxsD6KNE1SGUnOsEj04iunZJdsMKE9dpGd4muPuD8YgE2zuIrHWbu0AdOgjK
r+l9b53vZiyTre+ikiUUI7qXyJBh5cG2E9jXT6AfG4bT9xRhqN+jxFUhIBMOOXsqi2OODSI9hLGk
PetVAIPUvnStv05HX7vqJFMTNLwUohK7cyW8hu+w4MS9G4xC/U3U3VfiT1Xt9wbKah05y/kI/+be
VRvdAib8X9TGn5Sx6uj6zmiB2/vpMS+hu6IoUBrYX5Zxh3KsE4smSA5KJ34lZ2s2QJ+L4VEGEw/T
PGtwOeFh1C0nauacavxwhGK8graEOmqYU2mOHTatvU4o5dOxUq65C4j/6/6UXIUxJfVQPvJQu9XP
FfkaUc6RJshSolP6DwqCcTTOH+ZA2Dg9bD9fN/ieLU2FrsYbmD30LZj8MFPb3YjV3A3IeHzHIJ2r
D3FC8a5a2qjKEUXEzbd5hRy6pnq4mnGq8akLLYZonbnOJfanhPqE9x1WbNvD6HfNlLYh4ohT2KGc
QCz/Y5bAjtQsSdDVHs0OFqGx/lC2dyajjPsZEt4vfgefqz54kyy+3R5aMgq7vKUpklL8gnAtR6ca
oty8hSBeqsJnepqfeL4zcWP9nmILjReVYBcBPc3w9Dhn01qR6FtQUMHLfZYS+/xnmXnDMYePCxFX
ROIw2/mE6z8IPLeeC7/pz1HrnoCBLWBCTfUc3Gyd/uYhyqp4Nhgh3J1lhd9U4Isd39O8V12VgYa5
RvJ8dfKGC2rej87lmEyUW/hIpZVGYKhlX0FVugLNeZ9aobxJ7U0+dl4Qkq9E+W5bUk7Dzp9JJefm
DkNCE3mw6JNHsqpB9xjkBxDvrRivMVZUa8E4sEurfgKMvTKyvTeqZqTQuyyllLpg9PLZ6W3we1yB
C7SjG3KqsDMorGbRTj9upjbMQCTYB3qbcrHeccXHzr4svUyriLex0VEltTGdNqCDAvUQ5T5DjwX/
id5Dd+toDTSbM0wIv089QxNW6IXp3/tqqYqifzhbZX+OddiYDgjuIMRKBQQRJMtTBNOIDWD1+4tR
bg49vVDlaNVuJiLo9OxxDgzdIeN3UHCwlm0mytcmTFYkDO8nnJWfj5dPloenfY+amLsz3O03sOYf
PDMFdsT8tenfDZNEyKSXKj6ULf0ZTc0kK92vPkN7I5KB16ovfxBP5R74KR+8WT4izNypyS//280D
ZardPFGC/uJ/Lbo6nxXdOwb3JlCOrafE6PiCyXyXGUH4oFqe03ier8X8GDo7z1mcPaLzdNU1rpow
gkp1IM/ctcwdzgXaEUPjdA6UzcNcVqGWLGR1hxljbRzKshwhtvz8xVYUPfy5NOrPuTuaHCYZj6D4
LoB65WFAFRg73wJMDpWAG5Pr2qgfKSlYCR9cwlqKpkO2yidC6YppQiJkdkOJ+EQHJDwhdrW7zXPL
WrOiGD3r15K4i9pg6SJU4m21sLdP3HFL8hJU8sN2JoD/fJ4+ukPTM7TrUZlISyvrVoNT5B54c4mG
b3z6w7/bNt5LMSwjpSdN9GbTA5M3qtp+ne2UU0shSf8tS3izegYcPUfEUAdcwB+iwYBklJoQnBtZ
x9jLrhdQznie4DHzh88v/qFm4VqG+VQWY2njC74q7rBdEUoNVVZHeE30ADJhW14aVx2dUIAZsWvX
2CY1PCS6Ygsp8Zf1KDCyEQ7LBxHMX+kQ8pbbT59ZxIbohaOgibX/hwYI4zdhrSSkcye1Kzc/urup
z2RcCq/lqhzrOtLJ9TIoBjX96BqOHX6QbOUto/bswAjfBd3EWiL4HoUh5M4cLbv+mFbpmpuikdeC
RHEiJ55bFK2TkQCmACVT1yH62sUyMl/0vMGLtSOrot1fg7iCV9CAJMbQFBd9A/VAkxMX6rCtd+ZT
WiopXgtkNMsC0aUHSJt9nMBLSBJzZa6N/2p/UTiv69bRc3MtEJE/d9r41TkzpNkizsgO8RLEyV2T
Dowa3BDf2D1s82DY+iqF4SOO943W8NFFwgiD2B0RfFXeuFPMgXr6byNVAk2QASSPXSwy39xZtQm+
iL/auuW8Qp18PIs3luSRh7rkJ37m8Oe7kT+D2uLjHoifa/YU77tzIDuD+cP0MxtoTR6Rtrqbg2aS
LPvkpSQQF9byc8uUDRCTBSfEdJBNZ19bIg6dhN/IWYLU+zI7uv/JyxmrCwcWQGEunzcGlKngxlLE
vW/K4s7LvnoOvzgodfZBGMRm8e1piqg/r5kSWcYtRuKeXmmRnSrQ1oOjderCPE3gUQu9ulfgbOCN
KPH5zAlCS+kSOCtrp83lzFbtTz82kMBPqjVxFncD/0WKkGs3JSDiDj2CxE1vn9fkCGQDlzYxLMPc
DKBXBKkyQx6i1Q2f9IJqaZ6sz5Rc2cOikU0Yj5TI2dWv+GuXqM83TKkRBYHp84t9HSx3gL/xQ6G9
IofK3lHeuh44Tu4SRYsAy2we1RTzhean+r136i3AAc6Lmy6Jx6x7AiYsFQQhOWjyZ4xl83ZyHP47
POPmc8mzXr8pnjRnG6a8g6H2GelulqEyHjp/+FEkG5XNnMyoZBi0zIzgVvm3ht/xcQil0f3dbUPX
+WFfSKVJHqXmgrnxfyUleMpWsWKQhuc7kH6EV/W+cTR5Th/mCne/V8+79c/X0A2xg/qa+2AyFLEz
lmjcC74F+qfEImpvYRGv9WEo4+jWRfNsQBabtytWxx4n/gHEmXwMydoFPhqttFv10xWZyIWXVA29
DmRp20IWLGhqX3Sb+tziH5f7Ouzo2TBctSkfiWRqAjN7RPHSh171+dXe+6AWbAI8hQK1Udp8/jKZ
DU4aW+64mSxkBnm47tz9CEXnyj+EVd0OgMUk0aN8Yyl+Vb7GpCLafpMr2UZY27OhPPK4R763N1Qy
LLtUTMcqq0nOIG9b4TZLyFXqXF1KMDGhyyHtM5IX1S7qYh3Q+oESM9iar693XcbnMJYhX9Q3sNbq
WPJYK7NLZEwSA/8U9MHI9EX6M8f7L96oDdYMvSYSSJ8tWw8FTaV4S0DZI0tGNGQV/zEXpUWsCCiL
ayXwfYOYItEQsxx7mUFjVfhosAQ5A/JiuSnZUh0k7+OhzedFpM6ygN1KSgRl9Wz4L4W5NgCljpke
9A4nfR7xY5DlnF8ksLXsufpJVafhz63IjpoST+QnNhRtlIGZqyJkzI6c3PcNq1Mz70xd8QAvUbYP
78uw7KwFMIsspS0+IuyWVvW0RmeMh8FYd2+oGJ1xRJNgi+DO9VHxj9gQbTU5XTafgaY6oCIDVFS9
wWNdq+krOp5BFZIkxI+vX7k9i3qikQ+wOKreHQRWqsg9FdRMkq6uMXbDyJDjbKAX7TuELHYEVPGr
M3Hmpbf2h9B0jhl7bBoUOV7eHQWTmxArWU2a7rAB9ZiGC5AA9ir27UrBqWr0gTFnqUKBvvOTBcId
4Bl6ZiqoI7Cg6+8QhZZNJcgLEs495sgAhbOFpgywkoFNJUpkxedGhzXKNuf7kfDUY+ogbIQ1I20I
KbCimi4RM+95YGDx7OnxlYvqncWTCtw8/8wgyD/vwc1fBikfwQWEM3QXTcHistOdvPzntf5my/4D
w/CL6K+94GhasrumE+Ylfe3bF6VgR+nUCGgjgv77JwpARcwDByKMEYpSMtOgdYlL6dJtoORttMXZ
9laLg+HpvyT6O8WhhjIs/YgSNQxnz/ZxuDFz/nT7Eca3fQM/CLCDaSZPk0o71xhJE+uzhdES1pU4
ePYa3IdtqKqfGaN6TrsFqMVef7Sc7YZ1Z6OwTtpliW96xMTEnHW4iDoAo82NRrtjjWAGMuUHIpMJ
6Q7RPfOXXDHk/I90yL2lqXLSFomEpCFIsvjeyTSDfB/Uoy7LU01n16eQHUN3hnXmcQyL6ObwEYYo
HPs6bi8rl3HlCGZFC+RvFH7PnYODI7j2SkeCydXsJC4Y+Y6kwCO7Bg8zTC6Djkr9qrdKF23RC9YI
fl7jfoThQFf3+kETBp69RAX1M5Ttd1Zh+KlK29PHs+N5ytOje3oPGzc+plqekz1S8YvCok/0IzJy
/21T/Y8ll5ltwZqnqKoc2kR/ADra0NWhXJlY6Cj7iXzrjlmKQV3a2PEIC86CMrKBNUI1OUxxKzkP
RwfLKATFiKmHRqwTF+FKuv37AnyVXRJFvd/2yJyfmu2kA7RLc6PfiuPMcrwtulTaNzyqF7DAAuMV
7jfiVKjwL9LxZteVQK3alJyWjs45ARc7fVctun6K6jRBNDhEgqAk4BeKOzNgxsqKn7nQIqCCj09w
ohpqpaTqLAAae0fsRXY/iuUEa25/tlCWcnCBkR0UNo6uGV1YqqdqLxWCOnWVwXl0LDZhayTYGjwg
3IblbSt5GrED63FCjgLDueQzIUr9QBoa2CzzNptMu2SKKmOB6289A2PPedDYqC26l9Q3Tu0JjQqi
28cJBohoyF6urXWgy5kqUt0To63jV0jiqglytFOLlNqtvJ+N01dcMpKV72ra32hpDhqUqeSCZ6AV
inO5mYjTBeKV8rz6dhRgWQl79cUI0JUDxxcGsXbD4IiIGudAMlyRwWYowC4RxN4WPZQBGoaau3Hy
2H9DFElZyRRiBLa3N1HcJJ22RnQ6ZD0kAlu+KJSyIVbaUTHpe+3kvpbRQf0BBd5eLi+Pf/KxDAlt
bjYlxNjLhl3Fs7MS8ceiPQ9waJ7UKL646346wutK1DE9ov/ScsehUw1GX3vAUU8g5+Rzm7Qoxaxd
tiJqCvyfrGe0QVrytcalLbeaAvTYyxJI7GSbiW9U9awFVHfEnpYU2FrAua6d4eKhEnBXQevueFw/
WTu5oBp02ZD22r9iYZtPC1K8vNmIVs25Z8G5IavwrhprbsJZbjolnQIsXjpMqMkpCn0FXARixyu4
mjtrdyaAsfLPUvcxBvGO9hnDtwtvCC/IAvv/3TGjx1/U/ywWxRsHtDeB2+SJRe9VChPgi691DAi9
0SDzoK2L/LSf4c8ozwKuCCGdcW35RKSzDgEPMGU3/xqbHWXmyYfed9DvbxWJ7o5mcyb8vdQ8Wj+M
oLdyLwyrI7L4zB08dsHjXwg/eH0yMDvYnJRt7akvmYbvR2nKP8g5qN7cSi701SRYMr+DfQJNAGaq
cpY8ptZD/D74T8dwd3CtugDKgu7w1nr1WHGveZrVEFGcKNyYrJsAyMwL1xkTEMapOVckuFTD+i5l
3nZqU+wBJsS1WL9V+nl9M30Y9vCsdOHZ5faWmak0oEJofmAUmYve8RyBjGKooJ6rOfzdW7gOD1vq
9EcVMlXIDtH1dOpidmfIMyZmSSboermUAWAjHfgtiOs6XmDmKi/Y66R8dln7SdgmXXkJff/QYs2X
gZYnlagG4tOTYwnRxp6vsp/IBKyFhF5MNu4mBd5sS+HfOX2jbqKCuy+jvn7L8o85imEnVQtTSH2a
cISgVmkTAAgBklMRh2BCt/+GfxX+2HnMfHBUJfsOxtyS0w6V8phqCJ1OWXLIkAVIVC4GB+NMiPqI
1KeeC/kT67+9egEb8xxEE3sb2BQsyS4zc/r+Ijx9Y+k09QQtuN16/x+WnVKt4v1MT82yb6wGkK9B
/4K+T6ruD+Wuyi6Wo0RoZlOLKl/My0Y41VbYNSB2Xxzk9WwB9eVVkRSHqnr9rs22VhNJpEIr6Z8c
p9yQX8+HL4k6apQas7ht6QdNQrSSDRE0iJ+ocF938ufRvc7XhVSIBcMhJ3pFvcFYbUa+N+oOqFxI
0Fy6NlSkDE5bN1zjjFGY8H9x0YrFpNwraUa0B/d3FzQo6ZISIEL7zFCpjLyvZDpCObLvZMPy1nZw
t14jw/WJNhFVBMAT5IFbj5TH0RWXneKpWpuA9xckbtZDnHw4AahZHGzAiAIQzT2GoQ+YB91bC40j
B+Q8LLbeIGOajqOiJjcZhBqbUjM6nzly7H257mX85r9b3QDKM1oXjnndCWc+F7w1+iLk7HznX7IT
ncCCE51gzQIL9kw/iALBW+fL7BiYitR6KZLb9aFhnxkkq8YUNH7kOKl1K47cMpsaiCUu06MsIcgA
+1cHJ1QvUg/7ciLfUC+NvmWbCouYXSS+9ik3d+cgpXZa0A0eVFfcNUqDsjXMmTa2o41LJavlkQVL
/mLb7UMvhgMKO/N/zNORCOOMBvTzt5foPVZFEk4n4c5WvzoFufg0fRO7HXStTLJymyhmT/DXKvSK
PX/8sYB+OLxh32jXXjBn4W8LontfgCpWu5Cm93BvniAzkkf2PL1CVLvBdYJRa5DPo24lfDiv34//
66avn+gJP7FcMA1U61k9ux3ezRGPiUF+LZu7QiUmwyEgzR/HIP8Ko2jjHxbeovLCS9161KJrr0Um
vwqFgDmBN28CW17eIEOjLf/m5UTi6n7nsF7M/Mv+dM1jYwmpOPnzNgV5eqrOMhuTmqmg+5muj9QY
70AAIpDCknFw5Zq+KkzrrTQein2ThUlTPTKVoDycKTRe9LvTqFvtl6z6kvuDPiA3S5Xo6OO+vDwl
WKIe9xbXlvZkU2iry07M3ETcm8UFqI9AgtTLX8qtJip3zcVxj0I1QTncX2pOoV/p8Zdf8eYjX67D
kou8phlsCZvhwJMwGaex9tHLwKlt+8VfzIojHmoY9IcOa//ECEkcEn6O0YEFVtiGDhiC5YE1IEnc
K8OXt3fnBvGoG4wcadwMM9Umv1/YZduYR1zIY0Ud6iBNu2R7byVxcrp6iFIN+aOaIBJRFGqozX9R
Nt7XbahKeubd5IysRpHOLGezv0P0wJBy/YE6JVkIXqLMk/DmYaays2W3yXeZySojnwNM6LJD3pfs
ls5pTB5avfJCmzkwEh+HKEAJJTZEnhsHb5mMu3U3iAF1Stuqhqq8ZG41u2qjPwbjmE7xI+act0It
oOLbEbW9hvc3vLy6xvbCIO26GkuvC3QFBRiNa45BS6rw2N6hnTwTNVuLEPamJBxrhDLAm5GAG5i5
fW18wBEzZh3mXbLFvkwL6BPz9jLJp3K1aCEGmN2G08LpJkXGhhTUMKsnvrun3lFmrvVIrgqz3k50
2kXC2OeaaGIy6EMimoB0doRNUP4vTLGblgd98Sc1R15CP8me6tTQzbAUEDv9U/qv3N2XW3xDviaR
OyIQ2OyEBQ/Kq34ZyZhWS0V46pZqc/GfmSC0oyobXA4+zDIkG7H4TuonuVIzVE4gG9mQY/kL6VmG
SmViCM9ZZ8U1xdp36rM7WamxK9coF2UsiaH3YFlWpib/4+giGumwaQ1ch/h0y0kHoKdGF7U1XG5q
7iODwjotyr9PGnSccNWOe/zAmwYD7DuO5B0X0M1BlUbffLSFzDiyPxFUXF6+TbORiRT6u4my3P3N
tniagdHUjqAaoEUYUIIp8TkjYstOjotnVXrX5o+F6GW152aVCDDgeRBFD6UezJSQwzIpkqQOjUER
4JUfwwNs74zAz0P2mJacY5YpysbV5JF9oBJhv0l44h7Mzx8FT1LDPt+uIkK6lXx/3GuyLEd8ZIaq
uzc3Dr+/z1vDLinC2ifF2D86nI2Ip74LFelpJoOk3imMb56pRryowFq4KGJT6ei7K0pDDCm/Irzd
g6mzA7RvshAjq7aRUzQuUqkPUIkHQ2oeKBvEijuLwSohxCqpvdz3cxn1Ozws9/CuzzbOYiYSlLgm
FqFzXMORbQHSer8pQcdmXEWRgjSlmrd3+RgBsdbbjjITXTMjIDYXCVdRLxcgXHFDkxofZKWOwmKZ
sezOlJG0Ka+IMzbaoZ4B7Ao6Ek0GZBkeQFZUIvkC30w8FNHdiI9vBIjPxDSJ+xwP4Kx4K61UCbIl
KdUGlGKi/Mz5x2JfblYntjUlScTfd9tJ/CMZ7ZINR9ZIiC/s9yrRJ3MEaG+gGmjr86GGex0dPB6j
ifG7StLTG5s4Lf2XB1POBigCiF+yqsT2CPW6EezlxrC5PcT+w3XjxBIbb5z9vdgTaefwSabfnA1w
sZe60SWDMuqkyi2F54ozZVx2dgw+I19lj93BRLCwKM6gOZD2kR8BUCNeMkrPBNrcIuusMQTJQrs4
pMNXGtvc4yZxoBJ7TcRhN3Yw+He8Diok/vQ0q1s7wpKk3R3akIm6LFoXOcYAo4FaNDXeZp4MxXf7
G9xUmdaiOr6vGL97S/f1jE8hdmYgGAQSirADGA2dAMqM8BvmetPDb0iyUo9OhVFfVU+Wkm5r5OUq
q3xBHkctsXQISDUKg7Xy0rOzAE+CpHNg4ubwhgJqIpAbB1ZmeQOfkBOwujO0geGZX2wRTjNnsFhj
2OCh1WcsBBjxx1ImovbbY60zKezkd9s3EZosqqZujD5UEfVQjoTURYOY4OMHo8CQch4IUDmgut/y
P5T/mzVC5UcIx+DG9Xh9XGgZiHnu/lMJDoc9Muj7c/bW7o8B9xlPZ/E07k+zXGC4DK9k7+IDtNR4
7BORzsET2zSAqrTKRLLefKpkIL8ooXTqshluBQB5xUHl9+x+GWxUPV47q+QXx+y+C3IMrEw0ii4r
2kXDE5c40nLrbf0MbpPzRyBguMyHZdwm/qwtLQY28q8XbJ4XP4AXdYA5o8Mi2xnW58rOp2Zgikvr
IqAN4E79/m48e3EbVKuOvMrsX2pyT4UhGy9V5zwROKubmTrWQLyLrR86vxHFyMTm1El/KbEFsnPL
4QbQ5J0u3iuVlp7B4LXyFpPAWUXlf86n751sKNu57l9zy0b5s6U5NYmB4cUE4JVC7EYamteBvk+t
YAFToi89mTCxgOo2Iti8j9aiavMdukN5tlVMCZ5V95OwDyGkd1JsCsBetR5nmtu5PlXv6uvI9MQk
2Y82Fv6bueizNl7TNV39MjNZ2pYtmiKM9008gBjAe/HkVLsjDAIT63yCFFuHwjwqi/vNjvGk4MHj
k8118jLPwB1az0BVfuQJ5uQSV2HIwilm1MbVQvs/iIxNHBJWs4qsO5iakS75QkigaBSkHAMmUw6D
vHYyDelw7oTe1wWKTTdyxK5lZ4q/8zGxu8XROFMTZyZKeL3Jzjk1JNujmdLpQTBdIVwgSnW6YdeO
Y/wdDM6ilxMYO359suaw6iXnnwEN5C+1ZS0HZZ0EzZtKVRuoUrOWJUFfLPRQdEWXbEPhzgP3eK6r
LVsO6pbMm8wAQqC3j53VK7m7kXzHVgFKud7uwAXKtLPxknup/8z+RMOJuWNckrHtYMfv5wNc1gKx
80MQztH8bW4SFYwuoLPhqDz8oX/64UkuZxLHXo2XL3LyooIyRVrO9PPDzUUgh7C1Qn75JKqDH364
e/lJQjJsPYu9iFzYOo+lkChZL+m7c3Flo7e+89eeslhvD0mx7ZxwfnKV1XlSQWmAVEOfMtAHpnGR
ql+vgvqORU+jrblUkUG024jKblq6itxcGQ9KvhCoR7nysBdalbcf23nam2QML/2Vxr4twnefG8lO
09v+ibhbJ0LCsYdEtJCFWEtBwqK5uZumusWGiie2VFlVR+GsZk4HlWjyojVRzjxsXQ1r5qXg9kYV
MqRymFaIcIsgSnhXqz0dfWAaklsjH5lDB+X5Hp5cYQTqoexHZnuXXe5PYPTzN0XhvJxYMKrY8i63
rd3gNS1yMI2oLSO9fpT7EsLamI6d6hU6J0aRXUVpj74Czku72Ltg7gP4677K8a2P/eo34FpScKTH
0zuEndYsRvUkMN3zHuL6LOYGm+5xI6LJKgeb2duz2H5JFY+GMo9a8qxeh/KMztuCDIbUfDdCAYX6
yQDgQ/4PhDUvFOEC0TtHWMJ3kKDWZM56/50MZHtkjFQsT8tvRhlsIz3eXANgioMoh3GSL/2wboUm
jRTQbUF9CWJPdbel0vPyR/rfXpsyK7iTD5QJYQKGMpdBxmgj5+bf9D+g0H11765QlPkSH2SkcfTq
blK2Jbu+pAA6lk4AfF4ph2FqNZkF61WoGih9ScmdoxIeRK4if0WYOl5ogYZHL6F0lO87C/iWMDjr
FAV2d63cu8pGywOB45EOfTfZM/KjfvjCxMpe4uzJKCyjp9SDFFBONGzuc0FcFtrmVWFVsoaANd26
eeY/VePCuwRvAKmFgk+6ld4jYhXGRcSzQi9cJJfFSDIXc+nyyP9HBDKukLe8N9e6w/YCKbY3vSV4
VrpQDjR/LLz7LS+W29EzfLl/fpTZh4wE3LFr6oBEaMqFeMzuMxebm1VOrAiSLbbx80mCoWKCSsKL
Se9Jra9BnY0/BTpMWPr7ge//LPy/SRK3r7SydFPSpRMRHKYLaPtKx5aVtKNKmj7IsYLeOVdooaHM
7LkljdnPLlc21pUI/Rnvjct1NVzUDDo8qkd2PF970yBuziB9iZNY8S4A9gKgSC7o+/Bz/JAHMnuz
LcIZNr5WsPoWTU1xyctB05+dimDHzYZ+9pJff/in5lTW2YVxxibCkpdhthSv/MmWsv59CyCd0E5N
N+qfQ7eMcbhc6kBghALjo8sBOwLJF88WEePH9y8JQySPyYnh6F83y1MmsnCpCKAbHLQGRyx0KBLT
d4GkYammUItDwfv9B/ax7/9A8bddZgxTnIuPcfU5tc14OCK+hwB58ggu4XNcR1t2iHGm+AiZoPUH
jROpBsKXHt1w1N94yS/0SEVJSE6m7CYaJZRa6juTjU2cwbgR+yoE6+r94hHnq89wDjvbNP0qrL1v
luwEfXM0yn42B3BRilF7gvbwnUASC4k4qPU5nbMqjKkEjdyro8E3E8xm/Ba15OejVcklaY3tg1/W
q7nfrLaKLfiheFkZW/I7ZUuEiYb/bze6NX5ySEb7tdqPQCJzY2pgEgifJ4uPyF6gRTDZ4oCd3Iq6
Kz60JlhbK+MhKjr6GoxZvWRv2+3Hg108ZT750zRu6gqb/IZHcVGb1DPQsccFiPI4kZSbu3Q+7tKY
wMfC6XLFVgrrK0p79YzqcxsjP91Z44uFXGh9ZR9dnQB4Y7a1Jsh+czneRvQ637rTer2JY9QKP0E3
5zFVcO8A+T9Hd2k2bicSlztTtl7WQmwW+PZy4oxRqbKbWeQKbgltNs+8S7g/GXALFzXmTWD4OVcY
Wc4OCVszLUIhCdf9XjY36SDIhl9mPtV9eJPBjrWoNVa5f/bga4vf8iXS6mZWN/pWFbC5/TLHWhTg
+Fg5i7FPRmgnqh0wuMI7u2J8skfp/Af1uIJMQNDixTAmheLNWDqGB92TQ4COC9xQTJvHpxgaN3R0
K8SqneETVQsMepvgTfHyNSnjS6U60+z6vL9ZHVdeNo5DiDSw6Ve/ciiYHukMGJ3H4sKvyPO4EmWh
v64ZWyUNSWD6dCN3fq4V7OuIx9QF3V4FMAWtkKLHi9GmD43BxN1Wk8tnEKbwhzvjBx7ZY6O2Mz8p
nBuMX49NkmQ1li8NSDIN1dFmxWWSkVVilerWAuykpST1zc+kAKoB60FJ5BT2xGPBHwMxTWs0H8vR
TjIdQtM7s1bu7qZpHFUAFHU8QmTaMPdbT5DJiLHOftlW9LkBIjKW0TmAFlOyItNUrF38j5y92sZl
tXDvNpaeewFc8LiOLz9jlBKWMhmsqdAPm/PNNs074hz8VvqRwFye0ncU2gIAfG4V6HbzcYats4Q+
qEsC1VLwZH+eLrmoWN0xNfsDmhefGfcX4vHHzSsrrlha4190GcbP++kjc7jiM99PiPuuQbygV93E
fYmtddtx9gFATSWfJR9eNzcmX1Xl6JZ27KBTKWeOwGtyg21h6CmiNpVcbMmfRXqLFBY8mW6jYhya
nF0RHDVgzU+Hhwyy/MPxeRqyI1U4YtmisjiGDkh6cE+iVKhbouCAjXeBhTW3oV7cijH0HaS7XXra
jYAktbYLV9dACDM6h8mms9UvJ3Tkvqs97ze2s1V/+B3+/CGxcX7nfWLOhhpbP6TlTTOFQjye2SPB
6Q8dax3w6nULdnYP6ui0ja0ColEZETaKcQnRBp29/V/PiYJIhuFVpWYM4SjrqgF/bbrlI6fY43ry
IaThImeYtBitCGHxIFjMKqwszHZyR/3gMaq9SugsQ2l5ybw8HYjNYQRELVybDveL/VCb9F5I/lJ+
+ilCrt4us604eKrfhm6DfM1mZq4SkChtZHxj2RwzZxyTViACQGnoJDXWJbHmk0Zyt4oZUL+BnIvk
3ffGv/HwpaHku5WLsrrLEI05CqiDXN8IZxq0cmT2LiGZiezKT0obSlzHPPwR8yR5oeDnrIoJNKQ0
UPPm1r6ewoc1eDW/yJTWoMOJ86pCxkB8B3CRu5mIqttaliNgRylFcn6J331j8OeZzf/QuDWdqEz9
Agmn16HdpzxSAwPvyvzGeZZSqMV8BRX9plnq6+1Ok7RlXhN0INOwQ2oslpDDq21lubUNPcqoeFft
wCkEMk3vGaHkpq5+OYiGZX0eEFAv5nwDqjETwaVjb2W6iY/m5r4rsC2Qk09XZrrBUeOC5SOT8Xfp
PVFAkHBFOxE8HVGjoijnxEXLaX3glDk9iNrz0unecsG4HlKdvgE/yjLziYb0qCmrXVqYaqeWR1ut
lO/Ngd1WI9HfuPXsg8zDiKw8WgamIxTNSQbDPiOiYd3cjEdzL3WWTbQbpFXakkmjfmmfJhtY971R
1CVjA1NLLjIOqep6uZZAGRKrnbrVDefRgnPDXvbEH0fYNJOIzG4yHzUJDGcvVw4XhlqgJoCaOEMD
Qmj2WLmQ4z6Bnx+m11SzfexWImXi+B8FLRPeiAj/fDoLd1Wcr1DetCxsHl7vve/kmzI/noftXfWh
QA+TIhRRhCM+TZb6nWW/UVlobxg/ld9Y2Cl1DNXabR2s9q24nYoC8xUF+DBdpu+DeWeuZ39RDwom
vOPxkd8hULNc8Koy3zAHLsu0qkc8gtnUncWfYOJIivuSyoacu69+DCxasZjDbUfolSxOaGmHPh2e
mZ846pXAvwqbVVSJj6Dw+KfzEZDZMUzrGYPPeQJBssC8sFc0eR0oIKmUdahjQ4CPl0WjMwQA3nPg
oWaOXOPjJhRLoWICJfXAu5e7XuZWZZsObCDax7QztuMKioOQPX+SqXRf3k2VZFazfYXgNhrF+cPS
H3Fo6532mnNWQzeuy9d1/wugtyrLzvD1jykV6+qpYik+mgYm9PKkdEmThX0ojNXxIPhTLOq1t3vw
1M4J98SEnW/bWeHh9h4r100osbQft1pJ3nAClV3k539Z/h0y/yvbv1vocoO7GFbh2aqrgguLb1r2
yfQwgcLH/QRFAYDynFU/bO9CFT6/m4QVaDpJ+saSQgrgUKVl15v9vsGTnCKNOA2oNuaFln4nYb2h
Q9x/rBKds7IDMug6DzKtMEWpjKjKKT2l83giNjlXaaSvLsJA+wumOSeq7x1hahFAsmyPEd2MfKrz
ZXBpR9H41AkNKbSrSPiXM+p5qi+beuRBGuF4K5L3wP4oYN8WlFZVsY0xbTQvIRuyANC+fqKgNrwe
ivhkRa49pIhePeeHFG43kyi/A/0Zkx+VUoTTGgNsSwCBzj7D07PLecM0rDiscKewCNVuF2BtjmNa
WvGcfeFDtad8XbwDoZrl1Y7sPkrFLFc87kLXA4sV9H0iBFUn1aT0ImBy5B8mDtCHei7NL+t9Ny9j
RXJXuRjyAgt8coTWbd4oyECCZ4WtkL8qS0wQHMHZVWj4AqB0AksD8B4AhlAxxoRQ3YdbBj5TlQkj
F082lIEA6eDBBECaqinj+Rxv24S1Y9WTlUIdRNLrdnrJg81Z9/nYipXD3T4SEFWTsBPW0zHzZONd
38RJE0IC4sX/GYPhPtQgiMjOZEsoxaG1rIFz4GyDtkb6SkHT7/p4qtdwog7jqDSPQUmKX8oYfyU/
X2lvIXE5AdC2UIHB4j18b9Xo605YufL1gNgnxy9n5mZYVRBt94XST7AoCfY3Msh8hae7MfmB8CcW
4ahOBQf+DWhnxiUtIwrJvhuVYkahLg2/6ydBskteahcYXTlMt1QF87mUMRb25zzG5UyAPF22E0i1
I6sOD8YiXbA9Z8vgPHeBfq3ATEOStlJmU6hYVelhEERnoTnarMe2bGECJ1CsAVASzmYyu4aKwprB
n/ofRUkROIYiuVDYqwHgxg3siWXEjam378D/e23uLmChX1E3RlgF6Bg+2aLQDeop6YyXBEe08SvA
x0pSlUOdO4l5tFUDfE5H40VLmf31hkGEfx49msZuucp1UNNG18cFHKHClLQnkgmT7hXRma3KMIsS
LiJcivjviCC4+esAqjw7w+rUrRkr/sxErM39LciXIqcGGE/PTXHwHTzi7pZuEcy59m3Gs4958YLV
X54w1hJ5IJ3BItHaIeSuiIZjRJ68/Yh/7rSzSxHUlXVge+KfpD/laXX1X18+d7PEcPe2O3LS+YqR
2MLQK5kGHMq9Co6voBo+hiVJgFYBr1TmrcPkIAyGNMJsf3x3Jw+/S1RZwEhagDM9TSg2gXz/6yix
wFIQ5T8DMXIkukJTbA6uOWKQUjloGZ1eV37B1RFN3kmX+Uc/n7Wi1lOjeIlX397jFusY8ir3jr/3
uOkYzstY3hSHvjgyc/3WuCEZ8ihXB7zmYsPI+4xOBRT2n+fM0s6tndoJt5ZZIzFd9snQc0YfI7sj
InxX/dtza0MLAluzHpcHjHa2DjM26oFxTPu7he/9xj/oos7kn2tM6mRXnATZBVAU8aAWJZtrNvq2
T3dkHQhNpOIY/Ix2a5bw93qz57X+pMEYXFcAud4uJIYpmry6hvUA9mJjFbSoRR8SqFvu2JtPeOL/
CSVtmT78n5WhX8NKOUB8hyLoxDF/xtNrmThJOMJRZirJXJdNlDkx1ig0y8eZlqk3l1nm3qFHHCsv
2ZgSecbkiGOmtKawy/mIbSh7vNrKJr7epM1Oo/oH4pLRFeuSSzk/jMtF7+MQnDz19a+U69Agtl9w
rWjFdmlTrZS+ZadUJ4WJjsna3KpYbIGLO27K1/Px3qTM0Ni6tv7AjQOcniDfd9Rf1tXc8Azm3JFb
tjCBp7Tat1Q0rMyV25vmhZWsFcrKE7+2ZlqjFzdSYU8Rn3sduP5lanyT73ej0l3HjeXRvfa03APA
ytb7uxNVxUOJJiUSyE/u2gjX2UELlj5I9ASpQRDu186qk8Uk70nAG7AiJ3sMFhkeSqk599Lf/ebF
pOK9T1RsIKRBd39ERlc0RjO3IbBTk6WRgx3L0j9waFazRBBNwTLF1nXdh8GzFfpGRZhilp/q2vSx
7ERto5jAH6fiP6LuXXNQrDjmAgP8xxQH+wkHAibAzD1rB/oTG1U1kcCwGyxqgjv9AOpwtLLoslev
bBkezQn+4H6QX2nh9JsU9+vYhesLw2LDTbn96nKwlIfLK004JayZvLkaYyk1thcat6/9XDqASaOc
u09wKqNPAMrPOgLSNgWTCr3jHLeXMR2EyZo0yGXF9LFWfER2q4/HuOMLi5eEaRNVvjJkxZt240Cz
mlWXWB94kH0qBio0tja8mgg80/8u/RzrZGVR1fU3CWEX7pK9RogPubG6h5ojDELhkFYR7l1/aZ2q
hPKEIaR2C8rtGReBEpddjDEDd9J55+N3OB7KrbCZipWI4t1HwWhMmlnJIpixM8Ex5oNVt0DIefPx
7A6DtLOHrmx/BUe4rLLmbmOyj2Kr3fsNkrn/SApQ0rgFtlvJEABqIV5eqpJl0O8rNcruh2mSMsP2
XIM71sO0Z86d6xQuIzm1IMG6foBNHoVr4bF2TwJd0MMJLeH/243lk832SCfFyvAobi9a4hJTYtUQ
Tve2Xy6c7QUftfq7EEAdqm802BLHuzWKLjU1lhstHTj2MZGywG3iq9anRhqLywooBhWTH+eD2Nrf
yLror04gPakCW9thwwtzBa5cLED7OzMgq9EYgCeoaGJ345HnRJ0lHLHpGImNsSHWq038EPwO3H+b
VEpKGDi16M/vXKYSF4XcBITRMx62NsMG1+YF5BmfBmNq+t/aFPcHYgT6RPHVPEquw5wJmfu4qdX9
H2gMTkEt9tzCo2w384rYFZtyUwYIhWp8td8bT6Znd3/sic3k1FxU9hgA7JWH/eFPBJjmRos2MCrZ
JZguUfgxDEyYvUIi9F/pLN4dhNgaCg8Aup7aRVLy7uiroI8MYIAkGVcFnouee27LEn75nmFdcP3j
lYqJpEkXsoYnFNoVbvVwj6PsZKh3SEkQOwlzrFnUMAvvC0qS4XSAMYxEh7z+SMs0YMtEUp1ncG9z
1qruGMoyko9gS86qnnO5WbE7KIl5QuyFu365nddoDgPYji0zTXdH/OQn9V7kpL+mhqZT5xIktcmQ
w4PlMBX7jcQNWAo6toJhEC2L/E1+sdKofXM37tVDwRCFdtxkkOHOHNVnANRnxrKRwoQXLvdG0/w0
7Vaf54QHaH0nKYIPRD1tiVCJe51fxyzg8QGZxVm1xkU5t56nOSSxhl1nnEcv6PS7ICKggNpqYbTX
8spT69Udkykkv/4fcSCsnKX30U5Iyt52Jg3ILCA0EO9gD3vicQfaWQFyWBJRLI7T8APD3TIbkrt5
IIVo9oS51xq0A1rHRagpAaeIjGyef55u+LT3o9YnPGNwrfwAxSzUE2KjNIbIRdBDkyC1CwL4sdlz
X9AOzINIGwJpGKSAermncOZfrOrHNZq6xmT4xsmsyY47kjUrxB8VoeZxE+5oLxGg10bCpG17xhNv
bIWcVaVuIdz1QXmmazo0wMkZ3Vu8n3Ptz8W3eHJPpt4H9mftcfo10vUMPGORyuHRbw+yZVtVZx6Q
u+I0pPnUuQvMcVc0a0KGMXhcSFk7RSzcmfnjHCyeREuApga/KZJCahyW6Z5pBF3djAVLKJH8nBXb
g4DzibwStFQOyJdJLVH5Amjz01G28wyfJLFo7aojFANYe/Z7mK4f5DTF/ZS7Ed0KawI80/fz91RN
0PjXh/jo78rS4QdJ2NCLkQfxhcv7YSc1Lv8tiocvn+RUTeERSejn+kSrMApVfaA4UhTwvPll3wcM
AUk8WDK1fnA3/Kx33zmyzfmq17Ymz1dj52EeNQhk7fVVZHC9bG6GdHXU+kJqlnmp5frlYx0GK71m
wmMPxPthbNZ4TIAzh9cBNCaZdrSnX90R+3QOKTX3mU1hNQPCESmSPXDMGd/ecNAZi+jlP3OVMcrR
vGiC3Tp7Xj2dgdMD7N25y/0hDHHERZ1nS7JcpyCLuh3uJMi+bjBiRp8Npb91oTjeoQDqlzQZkpPb
nnlY0OeFU2rwmj7Cx4M3jWTsAunA2U8v7wpBqQQnUGc20LrnfysH3n160U7n3U6q/NC9BWip4wYB
FMpKRhw4bRUTXs8L/EXoatf69wQwKA+wCGzAQvV8WRzntZjbz8KxHhoFHkTuy1Gyf73QmQxk6bLK
96T/KpQPqU+ieMTIA8tBkSW+nLWkWIBA9kZQbURmaxo/2xaPO91SlFJB4f5AMDoyxF3wG+ULGWML
iowNKMKuexFeXM/dw1tOSmfqHvXS9eTyfQVxmN8NUYiQLKY9UGMPL8y30whLOD4WST5piRDTE1zs
fx4OQo8gPruWpizNCpCOAEGMAbxiTBaC8ultlI9XG6sd4+E9oIpREFi4pvH85sw4zcRO+ZX+YDuS
nEdr3Tp/hiQ3rZF2HxNqFVkmZExdZiSEk+UiqDxhuiFatleDktV/vOimivB6UDZxaE6XelDeksMP
vGbSI4wETt+8esqmyYJzCnb+gkJcGxXO+x0KsAmllS4Su3X7iGWaVAq/TCLSfZkzQYORayMFy/H6
91IvsxJMMEDIZbAX9Q3mBFX4ENdqvAIDvuhQ2TdHwYjpWMBpI8lVsq+xuBGnyHkz84Jpnw/dmGps
kjX3g9eeZU9n5zvJsZdhUPjSo5ojthzyNRVx9zJQV+EFDjZD/O3BD/k2p0QZ/h4VRyb5F30d0JoR
9g0giJI1VUIRkLYJuZ0uHj2lm3UtyqGS/DrRiSEPOXnoPeOjTuoFIjmNl//T1FNlDwt5X32jI34e
JoAdp3Nmzcg4sRVjtio8X9D/Eiba8zFkVlTAnI8GCSuhHsCLVnk7NFWGQdiQwa76xmq+e4tp1GJH
lrmfIpHuaLFDmFRIrAn7Lcrv4BZymhNmqI54T1KhlwKpznarR3oKEwx2FoETgX2g/xNAPWsLmh8+
9CE48MGb7Wk43PNe7fKegHgXn+S0zEP3EoDIeLN7XkUkp9T22h1bhFg0TuLYIB/EamP70JU1u+en
UeAt2REq+nphhynB6BS8WmwmdvDwrG7e4AqRE4FWKo8XTfHvED5Ztq1lwayXihDew18kmDJduH/E
GhfBDWGHLHq9wfhbV+XJyS1Bqok9w9XAabqz2wTKcg/hiDdQ6KcBqjenaO4n5I/bPfQTvP1SmVaD
yZ+PHvNy7Od+LDRuiQOI5PSTUzIS0QjSXDaxODmTzfJkEa4hqDctOCpH0aLe6xU3P7w54UVCeEp6
D89ofXyxBNPu+FHOkVwTFcBrp+M61gFroW8drqO+jY8I/R/PQUHr5wH+FPLn+6ZH3EZk0fRueeQN
2+kLX+W5MuO3uL+FYMQzgaX48GkOea5GdEIDoY2m85PhyiCd4GNRffHDEmCYKsXDYvT7bbJe85oU
kwmBQPOZR7vw6jBWrnl+2FRFb+DxVdbXJl+HP/Kl9D/oEGBa/l8m2zd942nVpqlOdo/ANlDAiB0p
SuXGxNrLHckUgOe/YJEA/ks9nS6yvRzRt3MwyA2QTkzU4ZiezCzQhzaF+cAixO3+tXkj7bGSEguU
jEy+5K3544javSVBhG6+j1npfpe375RDwprGm1hl2dDqc6PxiB6GHMdEh0lnvec1qxnm+H4pQoN8
1hhPJJZL4DFK1yhCOlncG1joduMH//Cnn6Mjdx1xsuNSaEcYRiSQs0SX3cv5lTYvw/NDMYms+HOZ
b3P2jI6mWGzOFwA7jet0a/up28TAJsy3gxu8y4V7VT5VbO1L9PZ14oLuSuYbDbxTADJ5YrRB+RZ7
/HZ9+WM4wERBUHDRyjVBxwwlEvO1uRwURBC2ZuS+JF0TIrjvBzpz94zjyuo+gSDxwkVbQAzAytLl
rgcDp2y+BwTXZPdmiuhCkeRPAZt+1rOgJKNp7EMiCEtPVu9kfMG2xtMm5YdV5S1HH2/eTZ9HPQhG
OfeWLLnFYkAxHSoZvNqU/2u8JexvFz7i2uxR3wMBXrcC9/JUl7sn3c2YUWHcsSGWVb41MTFv91f0
0DWxvYSFFFoP29PI7JHYVoNqtEpGpI3Drf895MyYLRyAO1eAVpOeX1qtKIOmIdfVJNA7EkoHc35w
9U7h8WDl8PiCug0xek/PNW62Jz0jHIyJGLoXSgop6vKKEpb+gEvl00cts2ZmY/bLp1EimiD0s6n8
eYa7oox+cMELW2Kys8voH7NWMHgwR9mZ9XAVq0ijkoFCEWQ7W1BLRBq7dXuGm157n+XvtCG4a0a6
zGEMe/vagqCIcyQLX5zk3e+2RdjnbFFGomg2WYc2JunRUFclOeAv9n/Wu7mPab1DtEgOcHAlZ7rO
BINSqVgcOk2+qenMa0mYL+J9M0ENqXQyATF1+tSFN38vgqK8Wqx3eZCXze8mB5NtqHaMLGzb7+xU
UwqU1KHznuy5heVqD94+yAx1t39YE5fN6SAaTd8QkE33cnFnTKsakZVjNlV47+hyoIK6Nlc9kaIB
Kwl2RwcOVbHbB4+ZArCL0izNHzUusDbFMZjU3WUbpKi14o+TN67gr5l7CTLcqLw9YFxYHuosYL9d
embmPju7JprT+idKU0/ktRnq+tDrksZ5UsgLoXrK/tEgogb1SlpJp8iM/Lz3cxqmTHpKEZEnRf0U
IBshzyxZnKtqYhk6asG2/krQrsam6U9SHqLFcKBY6B4S5RG5H5MKOffJGyz2UMcHDxl5RBKssGEv
x0HaiJBZ1D6TAsvU6j8VG0YXBtbFf/+w7l1ccelh5I6fR4q8fZVuyg/FV/aCd77WWk8YI6sChZF5
JLic7PbY5XaFf5f6pMtG2CpndwJ5QZuQLgGgCBZxdGzqlc4t3uEZU+U/QhW1YRXihnU+ypum2zcx
p4rzV1ryAnLEYMPcTe/pf71W/XVTY1GysggWjpPKTlw3test5xO7ty7Rn2dtXi/vzVcsx1ROAwOj
/jzNpRqYvyyWiwvyO5J6Dg6wMIvpf/WGgPxtVswc4M//Y8W6iJfMNt4LgwIU8E+gtlIHifhS8bFy
TJiUYjuWOUmlZFtR3dRXEIWP5DghtT+zTCRKYY+fVod0r2QfEiLiPNwU7BybUnGtgLFRL3TU5ssT
+TK+1dOjJ5JfyBz84aUl+lP9AI4l8g0jC0Ke3OQqgxfgTxMj+tu5oLBffYa/yGTN/w4IujAllQBA
XdZjzxvHQci3XELLQO4pRPeCmpsSDZf8m8BazbeKxXpoNKioSILk0GzuLGMaoxjnperm/87mK8Cu
0dOxh4V7PkyEZunYdWfmr6WTHnkm3yI3kC6qURTy9Rm9u6Vq8HRP6xUHOuoGsKtoNiIfCbYdyU5V
sSgQY1nSq1VMxYcGzyrEVowXiMwEWeC0red++NBExd/TyRQoiQkqD3goYdrwHnV8QQd79Fn3CPHL
jdXRTdikP6n5Fidz8WY93Psl69VWdNjKBImBT6hI/zOlu44T53rT5tILQwQv2h6I2YfP4Z0CUKk/
f2OH54DgwURxVEtmm5xf84SxlYymyp9f0j9BwiwcashF90hyq+7E99WMC7BN7zgUeWSZ2osi8huk
UDgZlSDH3bluuB9OCrVTP3VYOQ9UVrGzl14PWP1Vy6Bl03g1zNvFFe7QfaBB2B2/pRD0s5EZApOI
YC3ybX1KYQjKGzFgqFsWnfUJcJJ/gXZsH1NUp2bbfSuzb8h8TInEhTql3IoJBJ9M3emc6hb2vsag
bjVgeYOgoyAhp9vpbRj/gKgkFoupnyQ5db3/IMYiuGVKzKnzBZb7OYQKQxrvq+yo+x2fnDmdDh/I
V7/R0PZ3e1YRZ+CuOcS/Sv0MGWaWw8ohcO5BRRNIr+kcdc6eXn72bsupEgmGjVwG4hl/Wqgam+mZ
vXNjZ6Ombce0POe4EGdfYRPdyyGPwcIOXHorJWg8Jw/IHMNVkysUwrQS7FSsLkI4sAhObYRTZxd/
CGQXOtitbJTPloJs0g==

`protect end_protected

